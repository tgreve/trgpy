
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-06-10T03:07:33PDT



Photometric Data for RG J105239.84+572509.1

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|I (Cousins)         | 22.45     |+/-0.05 |mag                 |3.79E+14|  2.67E-06|+/-1.26E-07|Jy|2004ApJ...616...71S|1 sigma|    7900   A         | Broad-band measurement|| Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
2|K_s_ (2MASS)        | 18.89     |+/-0.10 |mag                 |1.38E+14|  1.85E-05|+/-1.79E-06|Jy|2004ApJ...616...71S|1 sigma|    2.17   microns   | Broad-band measurement|| Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
3|24 microns (MIPS)   | 150.      |+/-30   |uJy                 |1.27E+13|150.0E-06 |+/-30.0E-06|Jy|2009ApJ...694.1517D|1 sigma uncertainty|     23.68 microns   | Broad-band measurement|12 37 11.89 +62 22 11.8 (J2000)| Flux integrated from map|                                        |From new raw data
4|70 microns (MIPS)   |           |<9.3    |mJy                 |4.20E+12|          |9.3E-03|Jy|2009ApJ...699.1610H|3sigma|     71.42 microns   | Broad-band measurement|221804.42 +002154.4 (J2000)| Flux in fixed aperture|                                        |From new raw data
3|250 microns (SPIRE) | 25.02     ||milliJy             |1.20E+12|  2.50E-02||Jy|2010MNRAS.409L..13C|no uncertainty reported|       250 microns   | Broad-band measurement|10 52 39.840 +57 25 09.12 (J2000)| From fitting to map|                                        |From reprocessed raw data
4|350 microns (SPIRE) | 23.09     ||milliJy             |8.57E+11|  2.31E-02||Jy|2010MNRAS.409L..13C|no uncertainty reported|       350 microns   | Broad-band measurement|10 52 39.840 +57 25 09.12 (J2000)| From fitting to map|                                        |From reprocessed raw data
5|500 microns (SPIRE) | 20.83     ||milliJy             |6.00E+11|  2.08E-02||Jy|2010MNRAS.409L..13C|no uncertainty reported|       500 microns   | Broad-band measurement|10 52 39.840 +57 25 09.12 (J2000)| From fitting to map| 
5|850 microns (SCUBA) | -1.0      |+/-1.4  |mJy                 |3.53E+11|-1.0E-03  |+/-1.40E-03|Jy|2004ApJ...614..671C|1 sigma|       850 microns   | Broad-band measurement|105239.84 +572509.1 (J2000)| Flux integrated from map|                                        |From new raw data
7|850 microns (SCUBA) | 1.7       ||milliJy             |3.53E+11|  1.70E-03||Jy|2010MNRAS.409L..13C|no uncertainty reported|       850 microns   | Broad-band measurement|10 52 39.840 +57 25 09.12 (J2000)| From fitting to map|                                        |From reprocessed raw data
6|850 microns (SCUBA) |           |<2.7    |mJy                 |3.53E+11|          |2.7E-03|Jy|2004ApJ...614..671C|3rms sigma|       850 microns   | Broad-band measurement|105239.84 +572509.1 (J2000)| Flux integrated from map|                                        |From new raw data
7|1200 microns (MAMBO)|           |<2.1    |mJy                 |2.50E+11|          |2.1E-03|Jy|2004MNRAS.354..779G|3sigma uncertainty|      1200 microns   | Broad-band measurement|16 36 55.9 +40 59 12 (J2000)| Flux integrated from map|S/N = 3.66                              |From new raw data
8|1.4 GHz (VLA)       | 25.6      |+/-6.2  |microJy             |1.40E+09| 25.6E-06 |+/-6.2E-06|Jy|2006MNRAS.371..963B|1 sigma|       1.4 GHz       | Broad-band measurement|16 36 55.767 +40 59 09.97 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
