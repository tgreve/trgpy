
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-07-10T12:55:45PDT



Photometric Data for LEDA 2830476

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|H{beta} (VLT)       | 1.3E-15   ||erg/s/cm^2^         |6.17E+14|  1.30E+08||Jy-Hz|2011A&A...525A..43N|no uncertainty reported|      4861 A         | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|Broad line                              |From new raw data
2|H{alpha} (VLT)      | 5.5E-15   ||erg/s/cm^2^         |4.57E+14|  5.50E+08||Jy-Hz|2011A&A...525A..43N|no uncertainty reported|      6563 A         | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|Broad line                              |From new raw data
3|3.6 microns (IRAC)  | 68.4      |+/-7.1  | microJy            |8.44E+13|  6.84E-05|+/-7.10E-06|Jy|2007ApJS..171..353S|uncertainty|   3.550   microns   | Broad-band measurement|20 27 59.5 -21 40 56.90 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
4|4.5 microns (IRAC)  | 77.1      |+/-8.0  | microJy            |6.67E+13|  7.71E-05|+/-8.00E-06|Jy|2007ApJS..171..353S|uncertainty|   4.493   microns   | Broad-band measurement|20 27 59.5 -21 40 56.90 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
5|5.8 microns (IRAC)  | 86.8      |+/-10.9 | microJy            |5.23E+13|  8.68E-05|+/-1.09E-05|Jy|2007ApJS..171..353S|uncertainty|   5.731   microns   | Broad-band measurement|20 27 59.5 -21 40 56.90 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
6|8.0 microns (IRAC)  | 126.8     |+/-12.9 | microJy            |3.81E+13|  1.27E-04|+/-1.29E-05|Jy|2007ApJS..171..353S|uncertainty|   7.872   microns   | Broad-band measurement|20 27 59.5 -21 40 56.90 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
7|16 microns (IRS)    | 190.0     |+/-50.2 | microJy            |1.87E+13|  1.90E-04|+/-5.02E-05|Jy|2007ApJS..171..353S|uncertainty|      16   microns   | Broad-band measurement|20 27 59.5 -21 40 56.90 (J2000)| Flux in fixed aperture|6" diameter aperture                    |From reprocessed raw data
8|4.85 GHz            | 104       |+/-12   |milliJy             |4.85E+09|  1.04E-01|+/-1.20E-02|Jy|1994ApJS...90..179G|rms noise|4.85       GHz       | Broad-band measurement|202759.7 -214053 (J2000)| Modelled datum|                                        |From new raw data; Corrected for contaminating sources
9|1.4GHz (VLA)        | 342.2     |+/-10.3 |milliJy             |1.40E+09|  3.42E-01|+/-1.03E-02|Jy|1998AJ....115.1693C|uncertainty|    1.40   GHz       | Broad-band measurement|20 27 59.48 -21 40 57.0 (J2000)| Flux integrated from map|High Integral                           |From new raw data
10|408 MHz             | 1.28      |+/-0.08 |Jy                  |4.08E+08|  1.28E+00|+/-8.00E-02|Jy|1981MNRAS.194..693L|rms noise|408        MHz       | Broad-band measurement|202504.3 -215053 (B1950)| Modelled datum|                                        |From new raw data; Corrected for contaminating sources
11|365 MHz (Texas)     | 1.330     |+/-0.041|Jy                  |3.65E+08|  1.33E+00|+/-4.10E-02|Jy|1996AJ....111.1945D|internal error|365        MHz       | Broad-band measurement; obtained by interpolation over frequency|202504.204 -215055.29 (B1950)| Integrated from scans|Model:P;MFlag:+;EFlag:W;LFlag:+.        |From new raw data
