
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-06-16T16:22:30PDT



Photometric Data for DEEP2 13017707

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|K_s (Keck)          | 18.66     || mag                |1.39E+14|  2.13E-05||Jy|2007MNRAS.382..109T|no uncertainty reported|      2.15 microns   | Broad-band measurement|215.05412 +52.92598 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
2|24 microns (MIPS)   | 948       ||microJy             |1.27E+13|  9.48E-04||Jy|2010ApJ...719.1393D|no uncertainty reported|     23.68 microns   | Broad-band measurement|14 20 13.0 +52 55 33.3 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
