
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-03-28T04:01:20PDT



Photometric Data for COSMOS_J100054+023436,z=4.547

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
2|150              |   |<0.6     | uJy  | 2.00E15|  | 0.6E-6      |Jy |2003MNRAS.343..293M|1sigma uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
3|250              |   |<0.27     | uJy  | 1.20E15| | 0.09E-6      |Jy |2003MNRAS.343..293M|1sigma uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
4|380              |   |<0.03     | uJy  | 7.89E14| | 0.01E-6      |Jy |2003MNRAS.343..293M|1sigma uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
5|427              |   |<0.06     | uJy  | 7.03E14| | 0.02E-6      |Jy |2003MNRAS.343..293M|1sigma uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
6|446              |   |<0.03     | uJy  | 6.73E14| | 0.01E-6      |Jy |2003MNRAS.343..293M|1sigma uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
7|464              | 0.04  |+/-0.04| uJy  | 6.47E14| 0.04E-6| 0.04E-6 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
8|478              | 0.03  |+/-0.02| uJy  | 6.28E14| 0.03E-6| 0.02E-6 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
9|484              | 0.04  |+/-0.04| uJy  | 6.20E14| 0.04E-6| 0.04E-6 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
10|505              | 0.09  |+/-0.05| uJy  | 5.94E14| 0.09E-6| 0.05E-6 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
11|527              | 0.08  |+/-0.04| uJy  | 5.69E14| 0.08E-6| 0.04E-6 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
12|548              | 0.15  |+/-0.02| uJy  | 5.47E14| 0.15E-6| 0.02E-6 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
13|574              | 0.18  |+/-0.05| uJy  | 5.23E14| 0.18E-6| 0.05E-6 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
14|624              | 0.25  |+/-0.06| uJy  | 4.81E14| 0.25E-6| 0.06E-6 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
15|630              | 0.50  |+/-0.03| uJy  | 4.76E14| 0.50E-6| 0.03E-6 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
16|679              | 1.24  |+/-0.06| uJy  | 4.42E14| 1.24E-6| 0.06E-6 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
17|709nm            | 1.30  |+/-0.07| uJy  | 4.23E14| 1.30E-6| 0.07E-6 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
18|711nm            | 1.32  |+/-0.13| uJy  | 4.21E14| 1.32E-6| 0.13E-6 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
19|738nm            | 1.59  |+/-0.09| uJy  | 4.07E14| 1.59E-6| 0.09E-6 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
20|764nm            | 1.60  |+/-0.05| uJy  | 3.93E14| 1.60E-6| 0.05E-6 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
21|767nm            | 1.59  |+/-0.09| uJy  | 3.91E14| 1.59E-6| 0.09E-6 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
22|815nm            | 1.60  |+/-0.09| uJy  | 3.68E14| 1.60E-6| 0.09E-6 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
23|827nm            | 1.48  |+/-0.09| uJy  | 3.63E14| 1.48E-6| 0.09E-6 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
24|904nm            | 1.82  |+/-0.1| uJy  | 3.32E14| 1.82E-6| 0.1E-6 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
25|1.25um (Spitzer) | 2.4  |+/-0.8| uJy  | 2.40E14| 2.4E-6| 0.8E-6 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
26|2.15um (Spitzer) | 3.7  |+/-0.5| uJy  | 1.40E14| 3.7E-6| 0.5E-6 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
27|3.6um (Spitzer)  | 7.9  |+/-0.2| uJy  | 8.33E13| 7.9E-6| 0.2E-6 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
28|4.5um (Spitzer)  | 5.8  |+/-0.4| uJy  | 6.67E13| 5.8E-6| 0.4E-6 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
29|5.8um (Spitzer)  | 3.4  |+/-1.3| uJy  | 5.17E13| 3.4E-6| 1.3E-6 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
30|8.0um (Spitzer)  | 10. |+/-3.6| uJy  | 3.75E13| 10.E-6| 3.6E-6 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
31|24um (Spitzer)*  | 26.0 |+/-13.| uJy  | 1.25E13| 26.0E-6| 13.E-6 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
32|1.1mm (AzTEC)  | 4.8 |+/-1.5| mJy  | 2.73E11| 4.8E-3| 1.5E-3 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
33|1.25mm (MAMBO2)    | 3.41 |+/-0.67| mJy  | 2.4E11| 3.41E-3| 0.67E-3 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
34|83.3GHz (PDBI)     | 0.17 |0.08| mJy  | 83.3E9| 0.17E-3| 0.08E-3 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
34|41.7GHz (VLA)     |  |<150.| uJy  | 41.7E9| | 150.E-6 |Jy |2003MNRAS.343..293M|1sigma uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
34|1.4GHz (VLA)     | 45. |+/-9.| uJy  | 1.4E9| 45.E-6| 9.E-6 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
