
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-04-04T08:09:43PDT



Photometric Data for SMM J13123+4239

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|R (SUBARU)          | 24.7      |+/-0.3  |mag                 |4.76E+14|  4.11E-07|+/-1.14E-07|Jy|2006ApJS..167..103F|rms uncertainty|    6300   A         | Broad-band measurement| | Flux in fixed aperture|3" radius aperture                      |From new raw data
2|H{alpha} (UKIRT)    | 1.9E-19   |+/-0.1E-19| W/m^2^             |4.57E+14|  4.16E-08|+/-2.19E-09|Jy|2004ApJ...617...64S|uncertainty|      6563 A         | Line measurement; flux integrated over line; lines measured in emission|131232.31 +423949.5 (J2000)| Flux integrated from map|                                        |From new raw data
3|I (Cousins)         | 23.48     |+/-0.09 |mag                 |3.79E+14|  1.03E-06|+/-8.94E-08|Jy|2004ApJ...616...71S|1 sigma|    7900   A         | Broad-band measurement| | Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
4|z (SUBARU)          | 24.1      |+/-0.5  |mag                 |3.26E+14|  5.02E-07|+/-2.31E-07|Jy|2006ApJS..167..103F|rms uncertainty|    9200   A         | Broad-band measurement| | Flux in fixed aperture|3" radius aperture                      |From new raw data
5|J (2MASS)           | 21.75     |+/-0.23 |mag                 |2.40E+14|  3.18E-06|+/-7.50E-07|Jy|2004ApJ...616...71S|1 sigma|    1.25   microns   | Broad-band measurement| | Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
6|F160W (HST) AB      | 22.85     |+/-0.09 |mag                 |1.87E+14|  2.63E-06|+/-2.18E-07|Jy|2010MNRAS.405..234S|uncertainty|      1.60 microns   | Broad-band measurement|13 12 32.31 +42 39 49.5 (J2000)| Flux in fixed aperture|                                        |From new raw data
7|K_s_ (2MASS)        | 19.61     |+/-0.12 |mag                 |1.38E+14|  9.55E-06|+/-1.12E-06|Jy|2004ApJ...616...71S|1 sigma|    2.17   microns   | Broad-band measurement| | Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
8|3.6 microns (IRAC)  | 27.6      |+/-2.9  |microJy             |8.44E+13|  2.76E-05|+/-2.90E-06|Jy|2009ApJ...699.1610H|uncertainty|     3.550 microns   | Broad-band measurement|13 12 32.31 +42 39 49.5 (J2000)| Flux in fixed aperture|                                        |From new raw data
9|4.5 microns (IRAC)  | 43.8      |+/-4.6  |microJy             |6.67E+13|  4.38E-05|+/-4.60E-06|Jy|2009ApJ...699.1610H|uncertainty|     4.493 microns   | Broad-band measurement|13 12 32.31 +42 39 49.5 (J2000)| Flux in fixed aperture|                                        |From new raw data
10|5.8 microns (IRAC)  | 78.5      |+/-9.2  |microJy             |5.23E+13|  7.85E-05|+/-9.20E-06|Jy|2009ApJ...699.1610H|uncertainty|     5.731 microns   | Broad-band measurement|13 12 32.31 +42 39 49.5 (J2000)| Flux in fixed aperture|                                        |From new raw data
11|8.0 microns (IRAC)  | 197.0     |+/-20.0 |microJy             |3.85E+13|  1.97E-04|+/-2.00E-05|Jy|2009ApJ...699.1610H|uncertainty|     7.782 microns   | Broad-band measurement|13 12 32.31 +42 39 49.5 (J2000)| Flux in fixed aperture|                                        |From new raw data
12|850 microns (SCUBA) | 4.7       |+/-1.1  |milliJy             |3.53E+11|  4.70E-03|+/-1.10E-03|Jy|2005ApJ...622..772C|uncertainty|     850   microns   | Broad-band measurement|131232.31 +423949.5 (J2000)| Flux integrated from map|                                        |From new raw data
13|CO(3-2) line (IRAM) | |<1.4       |Jy km s^-1^         |3.46E+11| |4.26E-07|Jy|2005MNRAS.359.1165G|3 sigma|  2.3115             | Line measurement; flux integrated over line; lines measured in emission|... ... (J2000)| Flux integrated from map|                                        |From new raw data
14|1.4 GHz (VLA)       | 97        |+/-09   |microJy             |1.40E+09|  9.70E-05|+/-9.00E-06|Jy|2006ApJS..167..103F|uncertainty|     1.4   GHz       | Broad-band measurement|13 12 32.308 +42 39 49.58 (J2000)| Flux integrated from map|Corrected to the sky; see paper         |From new raw data
