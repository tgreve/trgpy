
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-02-19T12:04:08PST

z=2.56530

Photometric Data for SMM J14009+0252

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|0.2-2.0 keV (ROSAT)  | 4.1850E-14|+/-31.5%|erg/s/cm^2^         |3.15E+17|  1.33E-08|+/-4.19E-09|Jy|2000WGA...C...0000W|mean error| 1.3       keV       | Broad-band measurement|140050.7 +025201. (J2000)| Flux integrated from map|                                        |From reprocessed raw data; NED frequency assigned tomid-point of band in keV
2|F850LP (HST)         |           |>26.50  | mag                |3.17E+14| |5.50E-08|Jy|2008A&A...477...55H|3 sigma|      9445 A         | Broad-band measurement|14 00 57.530 +02 52 49.34 (J2000)| Flux in fixed aperture|                                        |From new raw data
3|SZ (VLT)             | 24.08     |+/-0.26 | mag                |2.83E+14|  4.15E-07|+/-9.95E-08|Jy|2008A&A...477...55H|rms uncertainty|      1.06 microns   | Broad-band measurement|14 00 57.530 +02 52 49.34 (J2000)| Flux in fixed aperture|                                        |From new raw data
4|J (VLT)              |           |>24.40  | mag                |2.40E+14| |2.76E-07|Jy|2008A&A...477...55H|3 sigma|      1.25 microns   | Broad-band measurement|14 00 57.530 +02 52 49.34 (J2000)| Flux in fixed aperture|                                        |From new raw data
5|H (VLT)              | 21.78     |+/-0.06 | mag                |1.82E+14|  1.99E-06|+/-1.10E-07|Jy|2008A&A...477...55H|rms uncertainty|      1.65 microns   | Broad-band measurement|14 00 57.530 +02 52 49.34 (J2000)| Flux in fixed aperture|                                        |From new raw data
6|K_s (VLT)            | 20.45     |+/-0.02 | mag                |1.39E+14|  4.41E-06|+/-8.12E-08|Jy|2008A&A...477...55H|rms uncertainty|      2.16 microns   | Broad-band measurement|14 00 57.530 +02 52 49.34 (J2000)| Flux in fixed aperture|                                        |From new raw data
7|3.6 microns (IRAC)   | 14.4      |+/-0.2  | microJy            |8.44E+13|  1.44E-05|+/-2.00E-07|Jy|2008A&A...477...55H|rms uncertainty|     3.550 microns   | Broad-band measurement|14 00 57.530 +02 52 49.34 (J2000)| Flux in fixed aperture|2.4" radius aperture                    |From reprocessed raw data
8|4.5 microns (IRAC)   | 23.0      |+/-0.3  | microJy            |6.67E+13|  2.30E-05|+/-3.00E-07|Jy|2008A&A...477...55H|rms uncertainty|     4.493 microns   | Broad-band measurement|14 00 57.530 +02 52 49.34 (J2000)| Flux in fixed aperture|2.4" radius aperture                    |From reprocessed raw data
9|5.8 microns (IRAC)   | 37.6      |+/-1.5  | microJy            |5.23E+13|  3.76E-05|+/-1.50E-06|Jy|2008A&A...477...55H|rms uncertainty|     5.731 microns   | Broad-band measurement|14 00 57.530 +02 52 49.34 (J2000)| Flux in fixed aperture|2.4" radius aperture                    |From reprocessed raw data
10|8.0 microns (IRAC)  | 50.9      |+/-1.6  | microJy            |3.81E+13|  5.09E-05|+/-1.60E-06|Jy|2008A&A...477...55H|rms uncertainty|     7.872 microns   | Broad-band measurement|14 00 57.530 +02 52 49.34 (J2000)| Flux in fixed aperture|2.4" radius aperture                    |From reprocessed raw data
11|12 microns (IRAS)   |           |<140    |mJy                 |2.50E+13|          |1.40E-01|Jy|1999ApJ...519..610D|3rms uncertainty reported| 20        cm        | Broad-band measurement|164502.36 +462625.5 (J2000)| Not reported in paper|                                        |Averaged from previously published data
12|24 microns (MIPS)   | 320.0     |+/-11.0 | microJy            |1.27E+13|  3.20E-04|+/-1.10E-05|Jy|2008A&A...477...55H|rms uncertainty|     23.68 microns   | Broad-band measurement|14 00 57.530 +02 52 49.34 (J2000)| Flux in fixed aperture|6" radius aperture                      |From reprocessed raw data
13|25 microns (IRAS)   |           |<155    | mJy                |1.20E+13|          |1.55E-01|Jy|2008A&A...477...55H|3rms uncertainty|     23.68 microns   | Broad-band measurement|14 00 57.530 +02 52 49.34 (J2000)| Flux in fixed aperture|6" radius aperture                      |From reprocessed raw data
14|60 microns (IRAS)   |           |<330    |mJy                 |5.00E+12| |3.30E-01|Jy|2008A&A...477...55H|3rms uncertainty|     23.68 microns   | Broad-band measurement|14 00 57.530 +02 52 49.34 (J2000)| Flux in fixed aperture|6" radius aperture                      |From reprocessed raw data
15|100 microns (IRAS)  |           |<415    |mJy                 |3.00E+12| |4.15E-01|Jy|1999ApJ...519..610D|3rms uncertainty| 20        cm        | Broad-band measurement|164502.36 +462625.5 (J2000)| Not reported in paper|                                        |Averaged from previously published data
16|450 microns (SCUBA) | 33        |        |milliJy             |6.66E+11|  3.30E-02| |Jy|2002MNRAS.331..495S|3rms uncertainty|     450   microns   | Broad-band measurement|140057.7 +025250 (J2000)| Flux integrated from map|                                        |From new raw data
17|450 microns (SCUBA) | 32.7      |+/-8.9  |milliJy             |6.66E+11|  3.27E-02|+/-8.9E-03|Jy|2002MNRAS.331..495S|uncertainty reported|     450   microns   | Broad-band measurement|140057.7 +025250 (J2000)| Flux integrated from map|                                        |From new raw data
18|450 microns (SCUBA) | -2        |+/-13   |milliJy             |6.66E+11| -2.00E-03|+/-1.30E-02|Jy|2007MNRAS.376.1073Z|uncertainty|     450   microns   | Broad-band measurement|14 00 57.5 +02 52 51 (J2000)| Flux integrated from map|                                        |From reprocessed raw data
19|850 microns (SCUBA) | 14.5      |        |milliJy             |3.53E+11|  1.45E-02| |Jy|2002MNRAS.331..495S|no uncertainty reported|     850   microns   | Broad-band measurement|140057.7 +025250 (J2000)| Flux integrated from map|                                        |From new raw data
20|850 microns (SCUBA) | 16.0      |        |milliJy             |3.53E+11|  1.60E-02| |Jy|2007MNRAS.376.1073Z|no uncertainty reported|     850   microns   | Broad-band measurement|14 00 57.5 +02 52 51 (J2000)| Flux integrated from map|S/N = 10.2                              |From reprocessed raw data
21|850 microns (SCUBA) | 15.6      |+/-1.9  |milliJy             |3.53E+11|  1.56E-02|+/-1.9E-03|Jy|2002MNRAS.331..495S|uncertainty reported|     850   microns   | Broad-band measurement|140057.7 +025250 (J2000)| Flux integrated from map|                                        |From new raw data
22|1350 microns (OVRO) | 5.57      |+/-1.72 |milliJy             |2.22E+11|  5.57E-03|+/-1.72E-03|Jy|2007MNRAS.376.1073Z|uncertainty reported|     850   microns   | Broad-band measurement|14 00 57.5 +02 52 51 (J2000)| Flux integrated from map|S/N = 10.2                              |From reprocessed raw data
18|146.5 GHz (IRAM)    | 10.2      |+/-1.3  |milliJy             |1.46E+11|  1.02E-02|+/-1.30E-03|Jy|2009ApJ...705L..45W|uncertainty|   146.469 GHz       | Broad-band measurement|| Flux integrated from map|                                        |From new raw data
20|87.9 GHz (IRAM)     | 5.4       |+/-0.9  |milliJy             |8.79E+10|  5.40E-03|+/-9.00E-04|Jy|2009ApJ...705L..45W|uncertainty|    87.888 GHz       | Broad-band measurement|| Flux integrated from map|                                        |From new raw data
23|32GHz (JVLA)        | 42.       |+/-20   |uJy                 |32.0E+9|  42.E-06|+/-20.E-06|Jy|2007MNRAS.376.1073Z|uncertainty reported|     850   microns   | Broad-band measurement|14 00 57.5 +02 52 51 (J2000)| Flux integrated from map|S/N = 10.2                              |From reprocessed raw data
24|1.05cm (OVRO)       |           |<0.54   |milliJy             |2.86E+10|  |0.54E-03 |Jy|2007MNRAS.376.1073Z|3rms uncertainty|     850   microns   | Broad-band measurement|14 00 57.5 +02 52 51 (J2000)| Flux integrated from map|S/N = 10.2                              |From reprocessed raw data
25|8GHz (JVLA)         | 91.       |+/-18   |uJy                 |8.00E+9|  91.E-06|+/-18.E-06|Jy|2007MNRAS.376.1073Z|uncertainty reported|     850   microns   | Broad-band measurement|14 00 57.5 +02 52 51 (J2000)| Flux integrated from map|S/N = 10.2                              |From reprocessed raw data
26|5GHz (JVLA)         | 151.      |+/-17   |uJy                 |5.00E+9|  151.E-06|+/-17.E-06|Jy|2007MNRAS.376.1073Z|uncertainty reported|     850   microns   | Broad-band measurement|14 00 57.5 +02 52 51 (J2000)| Flux integrated from map|S/N = 10.2                              |From reprocessed raw data
27|21.5cm (VLA)        | 529.      |+/-30   |uJy                 |1.40E+9|  529.E-06|+/-30.E-06|Jy|2007MNRAS.376.1073Z|uncertainty reported|     850   microns   | Broad-band measurement|14 00 57.5 +02 52 51 (J2000)| Flux integrated from map|S/N = 10.2                              |From reprocessed raw data
