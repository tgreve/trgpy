
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-07-10T12:50:32PDT



Photometric Data for LEDA 2826255

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|H{alpha} (VLT)      | 5.3E-15   ||erg/s/cm^2^         |4.57E+14|  5.30E+08||Jy-Hz|2011A&A...525A..43N|no uncertainty reported|      6563 A         | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|Broad line                              |From new raw data
2|3.6 microns (IRAC)  | 119.0     |+/-12.0 | microJy            |8.44E+13|  1.19E-04|+/-1.20E-05|Jy|2007ApJS..171..353S|uncertainty|   3.550   microns   | Broad-band measurement|10 19 49.0 -22 19 58.03 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
3|4.5 microns (IRAC)  | 179.0     |+/-18.0 | microJy            |6.67E+13|  1.79E-04|+/-1.80E-05|Jy|2007ApJS..171..353S|uncertainty|   4.493   microns   | Broad-band measurement|10 19 49.0 -22 19 58.03 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
4|5.8 microns (IRAC)  | 273.0     |+/-27.0 | microJy            |5.23E+13|  2.73E-04|+/-2.70E-05|Jy|2007ApJS..171..353S|uncertainty|   5.731   microns   | Broad-band measurement|10 19 49.0 -22 19 58.03 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
5|8.0 microns (IRAC)  | 360.0     |+/-36.0 | microJy            |3.81E+13|  3.60E-04|+/-3.60E-05|Jy|2007ApJS..171..353S|uncertainty|   7.872   microns   | Broad-band measurement|10 19 49.0 -22 19 58.03 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
6|20 GHz (ATCA)       | 57        |+/-4    |milliJy             |1.99E+10|  5.70E-02|+/-4.00E-03|Jy|2010MNRAS.402.2403M|rms uncertainty|    19.904 GHz       | Broad-band measurement|10 19 49.01 -22 19 59.3 (J2000)| Flux integrated from map|                                        |From new raw data
7|8 GHz (ATCA)        | 175       |+/-9    |milliJy             |8.00E+09|  1.75E-01|+/-9.00E-03|Jy|2010MNRAS.402.2403M|rms uncertainty|         8 GHz       | Broad-band measurement|10 19 49.01 -22 19 59.3 (J2000)| Flux integrated from map|                                        |From new raw data
8|5000 MHz            | 0.240     ||Jy                  |5.00E+09|  2.40E-01||Jy|1990PKS90.C...0000W|no uncertainty reported|    5000   MHz       | Broad-band measurement|10 17 27.8 -22 05 00 (B1950)| Integrated from scans|                                        |Homogenized from new and previously published data
9|5 GHz (ATCA)        | 305       |+/-15   |milliJy             |5.00E+09|  3.05E-01|+/-1.50E-02|Jy|2010MNRAS.402.2403M|rms uncertainty|         5 GHz       | Broad-band measurement|10 19 49.01 -22 19 59.3 (J2000)| Flux integrated from map|                                        |From new raw data
10|4.85 GHz            | 261       |+/-17   |milliJy             |4.85E+09|  2.61E-01|+/-1.70E-02|Jy|1994ApJS...90..179G|rms noise|4.85       GHz       | Broad-band measurement|101947.9 -221956 (J2000)| Modelled datum|                                        |From new raw data; Corrected for contaminating sources
11|2700 MHz            | 0.430     ||Jy                  |2.70E+09|  4.30E-01||Jy|1990PKS90.C...0000W|no uncertainty reported|    2700   MHz       | Broad-band measurement|10 17 27.8 -22 05 00 (B1950)| Integrated from scans|                                        |Homogenized from new and previously published data
12|1.4GHz (VLA)        | 673.2     |+/-20.2 |milliJy             |1.40E+09|  6.73E-01|+/-2.02E-02|Jy|1998AJ....115.1693C|uncertainty|    1.40   GHz       | Broad-band measurement|10 19 49.01 -22 19 59.8 (J2000)| Flux integrated from map|                                        |From new raw data
13|408 MHz             | 1.04      |+/-0.04 |Jy                  |4.08E+08|  1.04E+00|+/-4.00E-02|Jy|1981MNRAS.194..693L|rms noise|408        MHz       | Broad-band measurement|101727.1 -220453 (B1950)| Modelled datum|                                        |From new raw data; Corrected for contaminating sources
14|408 MHz             | 1.040     ||Jy                  |4.08E+08|  1.04E+00||Jy|1990PKS90.C...0000W|no uncertainty reported|     408   MHz       | Broad-band measurement|10 17 27.8 -22 05 00 (B1950)| Integrated from scans|                                        |Homogenized from new and previously published data
15|365 MHz (Texas)     | 0.993     |+/-0.028|Jy                  |3.65E+08|  9.93E-01|+/-2.80E-02|Jy|1996AJ....111.1945D|internal error|365        MHz       | Broad-band measurement; obtained by interpolation over frequency|101726.978 -220452.13 (B1950)| Integrated from scans|Model:P;MFlag:+;EFlag:+;LFlag:+.        |From new raw data
