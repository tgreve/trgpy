
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-05-27T08:12:11PDT



Photometric Data for GOODS J123629.13+621045.8

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|4.0-8 keV (Chandra) | 1.25E-15  | |ergs cm^-2^ s^-1^   |1.45E+18|  8.61E-11| |Jy|2003AJ....126..539A|no uncertainty reported|       6   keV       | Broad-band measurement|12 36 29.11 +62 10 45.9 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
2|4-8 keV (Chandra)   | 1.10E-15  |+/-4   %|erg cm^-2^ s^-1^    |1.45E+18|  7.59E-11|+/-3.03E-12|Jy|2001AJ....122.2810B|estimated error|       6   keV       | Broad-band measurement|12 36 29.11 +62 10 45.9 (J2000)| Flux in fixed aperture|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
3|2-10 keV (Chandra)  | 1.54E-15  | |erg/cm^2^/s         |1.45E+18|  1.06E-10| |Jy|2010MNRAS.401.2763L|no uncertainty reported|      6.00 keV       | Broad-band measurement|189.121180 62.179280 (J2000)| Modelled datum|                                        |From reprocessed raw data; NED frequency assigned tomid-point of band in keV
4|2-8 keV (Chandra)   | 2.22E-15  |+/-4   %|erg cm^-2^ s^-1^    |1.21E+18|  1.83E-10|+/-7.34E-12|Jy|2001AJ....122.2810B|estimated error|       5   keV       | Broad-band measurement|12 36 29.11 +62 10 45.9 (J2000)| Flux in fixed aperture|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
5|2.0-8 keV (Chandra) | 2.23E-15  | |ergs cm^-2^ s^-1^   |1.21E+18|  1.84E-10| |Jy|2003AJ....126..539A|no uncertainty reported|       5   keV       | Broad-band measurement|12 36 29.11 +62 10 45.9 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
6|0.5-8 keV (Chandra) | 2.31E-15  |+/-4   %|erg cm^-2^ s^-1^    |1.03E+18|  2.24E-10|+/-8.97E-12|Jy|2001AJ....122.2810B|estimated error|    4.25   keV       | Broad-band measurement|12 36 29.11 +62 10 45.9 (J2000)| Flux in fixed aperture|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
7|0.5-8 keV (Chandra) | 2.31E-15  | |ergs cm^-2^ s^-1^   |1.03E+18|  2.25E-10| |Jy|2003AJ....126..539A|no uncertainty reported|    4.25   keV       | Broad-band measurement|12 36 29.11 +62 10 45.9 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
8|2.0-4 keV (Chandra) | 0.70E-15  | |ergs cm^-2^ s^-1^   |7.25E+17|  9.65E-11| |Jy|2003AJ....126..539A|no uncertainty reported|       3   keV       | Broad-band measurement|12 36 29.11 +62 10 45.9 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
9|1.0-2 keV (Chandra) | 0.15E-15  | |ergs cm^-2^ s^-1^   |3.63E+17|  4.14E-11| |Jy|2003AJ....126..539A|no uncertainty reported|     1.5   keV       | Broad-band measurement|12 36 29.11 +62 10 45.9 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
10|0.5-2 keV (Chandra) | 0.17E-15  | |ergs cm^-2^ s^-1^   |3.02E+17|  5.62E-11| |Jy|2003AJ....126..539A|no uncertainty reported|    1.25   keV       | Broad-band measurement|12 36 29.11 +62 10 45.9 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
11|0.5-2 keV (Chandra) | 0.16E-15  |+/-4   %|erg cm^-2^ s^-1^    |3.02E+17|  5.30E-11|+/-2.12E-12|Jy|2001AJ....122.2810B|estimated error|    1.25   keV       | Broad-band measurement|12 36 29.11 +62 10 45.9 (J2000)| Flux in fixed aperture|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
12|0.5-1 keV (Chandra) | 0.03E-15  | |ergs cm^-2^ s^-1^   |1.81E+17|  1.65E-11| |Jy|2003AJ....126..539A|no uncertainty reported|    0.75   keV       | Broad-band measurement|12 36 29.11 +62 10 45.9 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
13|U (KPNO/MOSAIC) AB  | 26.11     |+/-0.25 |mag                 |8.44E+14|  1.31E-07|+/-3.01E-08|Jy|2005ApJ...635..853B|uncertainty|    3552   A         | Broad-band measurement|123629.13 +621045.8 (J2000)| Flux in fixed aperture|3" aperture                             |Averaged new and previously published data
14|U (KPNO) AB         | 26.1      | | mag                |8.22E+14|  1.32E-07| |Jy|2004AJ....127.3137C|no uncertainty reported| 3647.65   A         | Broad-band measurement|189.121490 +62.17957 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
15|F435W (HST) AB      | 21.957    |+/-0.018|mag                 |6.92E+14|  5.99E-06|+/-9.93E-08|Jy|2011ApJ...734..121S|uncertainty|      4333 A         | Broad-band measurement|189.121506 62.179565 (J2000)| Total flux|                                        |From reprocessed raw data
16|F435W (HST) AB      | 27.88     |+/-0.76 |mag                 |6.92E+14|  2.56E-08|+/-1.79E-08|Jy|2011ApJ...734..121S|uncertainty|      4333 A         | Broad-band measurement|189.121506 62.179565 (J2000)| Modelled datum|Central point source mag                |From reprocessed raw data
17|F435W (HST) AB      | 21.96     |+/-0.17 |mag                 |6.92E+14|  5.97E-06|+/-9.35E-07|Jy|2011ApJ...734..121S|uncertainty|      4333 A         | Broad-band measurement|189.121506 62.179565 (J2000)| Modelled datum|Host galaxy mag                         |From reprocessed raw data
18|B (SUBARU) AB       | 25.70     |+/-0.15 |mag                 |6.81E+14|  1.91E-07|+/-2.63E-08|Jy|2005ApJ...635..853B|uncertainty|    4400   A         | Broad-band measurement|123629.13 +621045.8 (J2000)| Flux in fixed aperture|3" aperture                             |Averaged new and previously published data
19|B (Subaru) AB       | 25.7      | | mag                |6.77E+14|  1.91E-07| |Jy|2004AJ....127.3137C|no uncertainty reported| 4427.60   A         | Broad-band measurement|189.121490 +62.17957 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
20|V (Subaru) AB       | 24.9      | | mag                |5.48E+14|  3.98E-07| |Jy|2004AJ....127.3137C|no uncertainty reported| 5471.22   A         | Broad-band measurement|189.121490 +62.17957 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
21|V (SUBARU) AB       | 24.98     |+/-0.09 |mag                 |5.42E+14|  3.70E-07|+/-3.07E-08|Jy|2005ApJ...635..853B|uncertainty|    5530   A         | Broad-band measurement|123629.13 +621045.8 (J2000)| Flux in fixed aperture|3" aperture                             |Averaged new and previously published data
22|R (SUBARU) AB       | 24.05     |+/-0.04 |mag                 |4.68E+14|  8.71E-07|+/-3.21E-08|Jy|2005ApJ...635..853B|uncertainty|    6400   A         | Broad-band measurement|123629.13 +621045.8 (J2000)| Flux in fixed aperture|3" aperture                             |Averaged new and previously published data
23|R (Keck II) AB      | 24.83     | | mag                |4.62E+14|  4.25E-07| |Jy|2004AJ....127.3121W|no uncertainty reported|   648.7   A         | Broad-band measurement|12 36 29.177 +62 10 46.06 (J2000)| Total flux|                                        |From new raw data
24|R (Subaru) AB       | 24.1      | | mag                |4.59E+14|  8.32E-07| |Jy|2004AJ....127.3137C|no uncertainty reported| 6534.16   A         | Broad-band measurement|189.121490 +62.17957 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
25|I (Cousins)         | 22.35     |+/-0.01 |mag                 |3.79E+14|  2.93E-06|+/-2.71E-08|Jy|2004ApJ...616...71S|1 sigma|    7900   A         | Broad-band measurement| | Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
26|I (SUBARU) AB       | 22.89     |+/-0.04 |mag                 |3.79E+14|  2.54E-06|+/-9.34E-08|Jy|2005ApJ...635..853B|uncertainty|    7900   A         | Broad-band measurement|123629.13 +621045.8 (J2000)| Flux in fixed aperture|3" aperture                             |Averaged new and previously published data
27|I (Subaru) AB       | 22.9      | | mag                |3.76E+14|  2.51E-06| |Jy|2004AJ....127.3137C|no uncertainty reported| 7975.89   A         | Broad-band measurement|189.121490 +62.17957 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
28|z' (Subaru) AB      | 22.4      | | mag                |3.31E+14|  3.98E-06| |Jy|2004AJ....127.3137C|no uncertainty reported| 9069.21   A         | Broad-band measurement|189.121490 +62.17957 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
29|z' (SUBARU) AB      | 22.36     |+/-0.04 |mag                 |3.30E+14|  4.13E-06|+/-1.52E-07|Jy|2005ApJ...635..853B|uncertainty|    9097   A         | Broad-band measurement|123629.13 +621045.8 (J2000)| Flux in fixed aperture|3" aperture                             |Averaged new and previously published data
30|J (Hale/WIRC) AB    | 21.39     |+/-0.05 |mag                 |2.40E+14|  1.01E-05|+/-4.65E-07|Jy|2005ApJ...635..853B|uncertainty|   1.250   microns   | Broad-band measurement|123629.13 +621045.8 (J2000)| Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
31|J (2MASS)           | 20.38     |+/-0.05 |mag                 |2.40E+14|  1.12E-05|+/-5.29E-07|Jy|2004ApJ...616...71S|1 sigma|    1.25   microns   | Broad-band measurement| | Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
32|F160W (HST) AB      | 21.23     |+/-0.03 |mag                 |1.87E+14|  1.17E-05|+/-3.23E-07|Jy|2010MNRAS.405..234S|uncertainty|      1.60 microns   | Broad-band measurement|12 36 29.13 +62 10 45.8 (J2000)| Flux in fixed aperture|                                        |From new raw data
33|HK' (UH) AB         | 20.5      | | mag                |1.58E+14|  2.29E-05| |Jy|2004AJ....127.3137C|no uncertainty reported|18947.38   A         | Broad-band measurement|189.121490 +62.17957 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
34|K_s (Hale/WIRC) AB  | 19.47     | |mag                 |1.39E+14|  5.92E-05| |Jy|2005ApJ...633..748R|no uncertainty reported|   2.150   microns   | Broad-band measurement|12 36 29.13 +62 10 45.8 (J2000)| Flux in fixed aperture|                                        |From new raw data
35|K_s_ (Hale/WIRC) AB | 19.93     |+/-0.02 |mag                 |1.39E+14|  3.87E-05|+/-7.13E-07|Jy|2005ApJ...635..853B|uncertainty|   2.150   microns   | Broad-band measurement|123629.13 +621045.8 (J2000)| Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
36|K_s_ (2MASS)        | 18.03     |+/-0.02 |mag                 |1.38E+14|  4.09E-05|+/-7.61E-07|Jy|2004ApJ...616...71S|1 sigma|    2.17   microns   | Broad-band measurement| | Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
37|3.6 microns (IRAC)  | 95.7      |+/-9.9  |microJy             |8.44E+13|  9.57E-05|+/-9.90E-06|Jy|2009ApJ...699.1610H|uncertainty|     3.550 microns   | Broad-band measurement|12 36 29.08 +62 10 45.7 (J2000)| Flux in fixed aperture|                                        |From new raw data
38|3.6 microns (IRAC)  | 98.14     | |microJy             |8.44E+13|  9.81E-05| |Jy|2010A&A...514A...9P|no uncertainty reported|     3.550 microns   | Broad-band measurement|189.121 62.180 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
39|3.6 microns (IRAC)  | 97.00     |+/-4.85 |microJy             |8.44E+13|  9.70E-05|+/-4.85E-06|Jy|2011AJ....141....1T|rms uncertainty|     3.550 microns   | Broad-band measurement|189.121307 62.179440 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
40|3.6 microns IRAC AB | 18.96     |+/-0.04 |mag                 |8.44E+13|  9.46E-05|+/-3.49E-06|Jy|2005ApJ...635..853B|uncertainty|   3.550   microns   | Broad-band measurement|123629.13 +621045.8 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged new and previously published data
41|N4 (AKARI)          | 84.08     | |microJy             |6.92E+13|  8.41E-05| |Jy|2010A&A...514A...9P|no uncertainty reported|      4.33 microns   | Broad-band measurement|189.121 62.180 (J2000)| Flux in fixed aperture|                                        |From new raw data
42|4.5 microns (IRAC)  | 89.4      |+/-9.2  |microJy             |6.67E+13|  8.94E-05|+/-9.20E-06|Jy|2009ApJ...699.1610H|uncertainty|     4.493 microns   | Broad-band measurement|12 36 29.08 +62 10 45.7 (J2000)| Flux in fixed aperture|                                        |From new raw data
43|4.5 microns (IRAC)  | 88.33     | |microJy             |6.67E+13|  8.83E-05| |Jy|2010A&A...514A...9P|no uncertainty reported|     4.493 microns   | Broad-band measurement|189.121 62.180 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
44|4.5 microns (IRAC)  | 86.80     |+/-4.34 |microJy             |6.67E+13|  8.68E-05|+/-4.34E-06|Jy|2011AJ....141....1T|rms uncertainty|     4.493 microns   | Broad-band measurement|189.121307 62.179440 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
45|4.5 microns IRAC AB | 19.02     |+/-0.04 |mag                 |6.67E+13|  8.95E-05|+/-3.30E-06|Jy|2005ApJ...635..853B|uncertainty|   4.493   microns   | Broad-band measurement|123629.13 +621045.8 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged new and previously published data
46|5.8 microns (IRAC)  | 77.9      |+/-7.9  |microJy             |5.23E+13|  7.79E-05|+/-7.90E-06|Jy|2009ApJ...699.1610H|uncertainty|     5.731 microns   | Broad-band measurement|12 36 29.08 +62 10 45.7 (J2000)| Flux in fixed aperture|                                        |From new raw data
47|5.8 microns (IRAC)  | 76.03     | |microJy             |5.23E+13|  7.60E-05| |Jy|2010A&A...514A...9P|no uncertainty reported|     5.731 microns   | Broad-band measurement|189.121 62.180 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
48|5.8 microns (IRAC)  | 76.00     |+/-3.82 |microJy             |5.23E+13|  7.60E-05|+/-3.82E-06|Jy|2011AJ....141....1T|rms uncertainty|     5.731 microns   | Broad-band measurement|189.121307 62.179440 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
49|5.8 microns IRAC AB | 19.21     |+/-0.10 |mag                 |5.23E+13|  7.52E-05|+/-6.92E-06|Jy|2005ApJ...635..853B|uncertainty|   5.731   microns   | Broad-band measurement|123629.13 +621045.8 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged new and previously published data
50|8.0 microns (IRAC)  | 74.1      |+/-7.7  |microJy             |3.85E+13|  7.41E-05|+/-7.70E-06|Jy|2009ApJ...699.1610H|uncertainty|     7.782 microns   | Broad-band measurement|12 36 29.08 +62 10 45.7 (J2000)| Flux in fixed aperture|                                        |From new raw data
51|8 microns (IRAC)    | 70.62     | |microJy             |3.81E+13|  7.06E-05| |Jy|2010A&A...514A...9P|no uncertainty reported|     7.872 microns   | Broad-band measurement|189.121 62.180 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
52|8.0 microns IRAC AB | 19.34     |+/-0.06 |mag                 |3.81E+13|  6.67E-05|+/-3.69E-06|Jy|2005ApJ...635..853B|uncertainty|   7.872   microns   | Broad-band measurement|123629.13 +621045.8 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged new and previously published data
53|8.0 microns (IRAC)  | 72.10     |+/-3.64 |microJy             |3.81E+13|  7.21E-05|+/-3.64E-06|Jy|2011AJ....141....1T|rms uncertainty|     7.872 microns   | Broad-band measurement|189.121307 62.179440 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
54|S11 (AKARI)         | 75.10     | |microJy             |2.87E+13|  7.51E-05| |Jy|2010A&A...514A...9P|no uncertainty reported|     10.45 microns   | Broad-band measurement|189.121 62.180 (J2000)| Flux in fixed aperture|                                        |From new raw data
55|11 microns (AKARI)  | 75.0      |+/-15   | microJy            |2.73E+13|  7.50E-05|+/-1.50E-05|Jy|2009MNRAS.394..375N|uncertainty|        11 microns   | Broad-band measurement|12 36 29.16 +62 10 46.46 (J2000)| Flux integrated from map|                                        |From new raw data
56|16 microns (IRS)    | 463.0     |+/-18.3 |microJy             |1.90E+13|  4.63E-04|+/-1.83E-05|Jy|2011AJ....141....1T|rms uncertainty|      15.8 microns   | Broad-band measurement|189.121307 62.179440 (J2000)| From fitting to map|                                        |From new raw data
57|16 microns (IRS)    | 465.00    | |microJy             |1.87E+13|  4.65E-04| |Jy|2010A&A...514A...9P|no uncertainty reported|        16 microns   | Broad-band measurement|189.121 62.180 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
58|16 microns (IRS)    | 465       |+/-25   | microJy            |1.87E+13|  4.65E-04|+/-2.50E-05|Jy|2009MNRAS.394..375N|uncertainty|        16 microns   | Broad-band measurement|12 36 29.16 +62 10 46.46 (J2000)| Flux integrated from map|                                        |Averaged from previously published data
59|18 microns (AKARI)  | 434       |+/-33   | microJy            |1.67E+13|  4.34E-04|+/-3.30E-05|Jy|2009MNRAS.394..375N|uncertainty|        18 microns   | Broad-band measurement|12 36 29.16 +62 10 46.46 (J2000)| Flux integrated from map|                                        |From new raw data
60|L18W (AKARI)        | 433.77    | |microJy             |1.63E+13|  4.34E-04| |Jy|2010A&A...514A...9P|no uncertainty reported|     18.39 microns   | Broad-band measurement|189.121 62.180 (J2000)| Flux in fixed aperture|                                        |From new raw data
61|24 microns (MIPS)   | 699.0     |+/-71.0 |microJy             |1.27E+13|  6.99E-04|+/-7.10E-05|Jy|2009ApJ...699.1610H|uncertainty|     23.68 microns   | Broad-band measurement|123629.13 +621045.8 (J2000)| Flux in fixed aperture|                                        |From new raw data
62|24 microns (MIPS)   | 720.49    | |microJy             |1.27E+13|  7.21E-04| |Jy|2010A&A...514A...9P|no uncertainty reported|     23.68 microns   | Broad-band measurement|189.121 62.180 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
63|24 microns (MIPS)   | 730.0     |+/-12.7 |microJy             |1.27E+13|  7.30E-04|+/-1.27E-05|Jy|2011AJ....141....1T|rms uncertainty|     23.68 microns   | Broad-band measurement|189.121307 62.179440 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
64|24 microns (Spitzer)| 724       |+/-12   |microJy             |1.27E+13|  7.24E-04|+/-1.20E-05|Jy|2011ApJ...726...93R|uncertainty|     23.68 microns   | Broad-band measurement|12 36 29.13 +62 10 45.8 (J2000)| Not reported in paper|                                        |Averaged from previously published data
65|70 microns (MIPS)   | |<1.8       |mJy             |4.20E+12| |1.80E-03|Jy|2009ApJ...699.1610H|3 sigma|     71.42 microns   | Broad-band measurement|123629.13 +621045.8 (J2000)| Flux in fixed aperture|                                        |From new raw data
66|850 microns (SCUBA) | 5.0       |+/-1.3  |milliJy             |3.53E+11|  5.00E-03|+/-1.30E-03|Jy|2005ApJ...622..772C|uncertainty|     850   microns   | Broad-band measurement|123629.13 +621045.8 (J2000)| Flux integrated from map|                                        |From new raw data
67|850 microns (SCUBA) | 4.6       |+/-1.2  |milliJy             |3.53E+11|  4.60E-03|+/-1.20E-03|Jy|2005MNRAS.358..149P|uncertainty|     850   microns   | Broad-band measurement|12 36 28.7 +62 10 47 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
68|1.4 GHz (VLA)       | 81        | |microJy             |1.40E+09|  8.10E-05| |Jy|2005MNRAS.358.1159M|no uncertainty reported|     1.4   GHz       | Broad-band measurement|12 36 29.1240 +62 10 45.984 (J2000)| Flux integrated from map|                                        |From new raw data
69|1.4 GHz (VLA)       | 91        |+/-13   | microJy            |1.40E+09|  9.10E-05|+/-1.30E-05|Jy|2006MNRAS.371..963B|1 sigma|       1.4 GHz       | Broad-band measurement|12 36 29.159 +62 10 45.83 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
70|1.4 GHz (VLA)       | 100.8     |+/-12.9 |microJy             |1.40E+09|  1.01E-04|+/-1.29E-05|Jy|2010ApJS..188..178M|uncertainty|       1.4 GHz       | Broad-band measurement|12 36 29.05 +62 10 45.8 (J2000)| Total flux; Beam filling or dilution corrected|Major=2.8"; Minor=1.0"; PA=75 deg       |From new raw data
71|1.4 GHz             | 81.4      |+/-8.7  |microJy             |1.40E+09|  8.14E-05|+/-8.70E-06|Jy|2000ApJ...533..611R|1 sigma|1.4        GHz       | Broad-band measurement; broad-band flux derived by integration over spectrum; synthetic band|123629.134 +621045.79 (J2000)| Flux integrated from map; Pointing and beam filling|                                        |From new raw data; Corrected for contaminating sources
