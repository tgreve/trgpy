
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-05-28T01:42:09PDT



Photometric Data for H-ATLAS J090311.6+003906

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|0.48 microns (INT)  | 26.0      |+/-0.3  |microJy             |6.25E+14|  2.60E-05|+/-3.00E-07|Jy|2011ApJ...732L..35C|uncertainty|      0.48 microns   | Broad-band measurement|10 57 51.1 +57 30 27 (J2000)| Flux in fixed aperture|                                        |From new raw data
2|0.63 microns (INT)  | 46.5      |+/-0.6  |microJy             |4.76E+14|  4.65E-05|+/-6.00E-07|Jy|2011ApJ...732L..35C|uncertainty|      0.63 microns   | Broad-band measurement|10 57 51.1 +57 30 27 (J2000)| Flux in fixed aperture|                                        |From new raw data
3|0.76 microns Subaru | 47.9      |+/-0.3  |microJy             |3.94E+14|  4.79E-05|+/-3.00E-07|Jy|2011ApJ...732L..35C|uncertainty|      0.76 microns   | Broad-band measurement|10 57 51.1 +57 30 27 (J2000)| Flux in fixed aperture|                                        |From new raw data
4|i (Subaru) AB       | 22.72     |+/-0.01 |mag                 |3.91E+14|  2.96E-06|+/-2.73E-08|Jy|2011ApJ...738..125G|uncertainty|   7671    A         | Broad-band measurement|| Modelled datum|                                        |From new raw data
5|2.2 microns (Keck)  | 63.1      |+/-2.0  |microJy             |1.36E+14|  6.31E-05|+/-2.00E-06|Jy|2011ApJ...732L..35C|uncertainty|       2.2 microns   | Broad-band measurement|10 57 51.1 +57 30 27 (J2000)| Flux in fixed aperture|                                        |From new raw data
1|4.5 microns (IRAC)  | 376.0    |+/-6.0   |microJy             |6.67E+13 | 376.0E-06  |+/-6.0E-06 |Jy |2011ApJ...728L...4H|uncertainty|     4.493 microns   | Broad-band measurement|09 03 11.6 +00 39 06 (J2000)| Flux in fixed aperture|                                        |From new raw data
2|5.8 microns (IRAC)  | 442.0    |+/-11.0  |microJy             |5.23E+13 | 442.0E-06  |+/-11.0E-06|Jy|2009AJ....137.3884R|uncertainty|     5.731 microns   | Broad-band measurement|249.244975 40.957682 (J2000)| Flux integrated from map|                                        |From new raw data
3|8.0 microns (IRAC)  | 558.0    |+/-16.0  |microJy             |3.85E+13 | 558.0E-06  |+/-16.0E-06|Jy|2009ApJ...699.1610H|uncertainty|     7.782 microns   | Broad-band measurement|16 36 58.75 +40 57 27.8 (J2000)| Flux in fixed aperture|                                        |From new raw data
4|MIPS 24 microns     | 5.5      |+/-0.4   |mJy                 |1.25E+13 |   5.5E-03  |+/-0.4E-03 |Jy|1990IRASF.C...0000M|3sigma uncertainty| 25        microns   | Broad-band measurement|115813.1 +302058 (B1950)| Flux in fixed aperture|                                        |From new raw data
5|70 microns (MIPS)   | 22.2     |+/-3.0   |mJy                 |4.20E+12 |  22.2E-03  |+/-3.0E-03 |Jy|2009A&A...502..541E|uncertainty reported|     71.42 microns   | Broad-band measurement| | Flux in fixed aperture|Tentative detection                     |From reprocessed raw data 
6|160 microns (MIPS)  | 310.0    |+/-8.0   |mJy                 |1.92E+12 | 310.0E-03  |+/-8.0E-03|Jy|2009A&A...502..541E|3 sigma|     155.9 microns   | Broad-band measurement| | Flux in fixed aperture|                                        |From reprocessed raw data
7|250 microns (SPIRE) | 425.0    |+/-10.0  |mJy                 |1.199e+12|  425.0E-03 |+/-10.0e-03|Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
8|350 microns (SPIRE) | 340.0    |+/-10.0  |mJy                 |8.565e+11|  340.0E-03 |+/-10.0e-03|Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
9|500 microns (SPIRE) | 233.0    |+/-11.0  |mJy                 |5.996e+11|  233.0E-03 |+/-11.0e-03|Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
10|880 microns (SMA)   | 52.8     |+/-0.5   |mJy                 |3.40E+11 |  52.8E-03  |+/-0.5E-03|Jy|2010ApJ...709..210K|uncertainty|      870  microns   | Broad-band measurement|16 35 55.67 +66 12 59.51 (J2000)| Flux integrated from map|                                        |From new raw data
11|1050 microns (Z-SPEC)| 27.5     |+/-0.6   |mJy                |2.86E+11 |  27.5E-03  |+/-0.6E-03|Jy|2010ApJ...709..210K|uncertainty|      870  microns   | Broad-band measurement|16 35 55.67 +66 12 59.51 (J2000)| Flux integrated from map|                                        |From new raw data
12|1150 microns (Z-SPEC)| 20.4     |+/-0.5   |mJy                |2.61E+11 |  20.4E-03  |+/-0.5E-03|Jy|2010ApJ...709..210K|uncertainty|      870  microns   | Broad-band measurement|16 35 55.67 +66 12 59.51 (J2000)| Flux integrated from map|                                        |From new raw data
13|1250 microns (Z-SPEC)| 16.2     |+/-0.5   |mJy                |2.40E+11 |  16.2E-03  |+/-0.5E-03|Jy|2010ApJ...709..210K|uncertainty|      870  microns   | Broad-band measurement|16 35 55.67 +66 12 59.51 (J2000)| Flux integrated from map|                                        |From new raw data
14|1350 microns (Z-SPEC)| 12.0     |+/-0.5   |mJy                |2.22E+11 |  12.0E-03  |+/-0.5E-03|Jy|2010ApJ...709..210K|uncertainty|      870  microns   | Broad-band measurement|16 35 55.67 +66 12 59.51 (J2000)| Flux integrated from map|                                        |From new raw data
15|1450 microns (Z-SPEC)| 9.9     |+/-0.5   |mJy                |2.07E+11 |  9.9E-03  |+/-0.5E-03|Jy|2010ApJ...709..210K|uncertainty|      870  microns   | Broad-band measurement|16 35 55.67 +66 12 59.51 (J2000)| Flux integrated from map|                                        |From new raw data
16|3400 microns (CARMA)| 0.61     |+/-0.19   |mJy                |8.82E+10 |  0.61E-03  |+/-0.19E-03|Jy|2010ApJ...709..210K|uncertainty|      870  microns   | Broad-band measurement|16 35 55.67 +66 12 59.51 (J2000)| Flux integrated from map|                                        |From new raw data
17|1.4 GHz (VLA)       | 1.8      |+/-0.7   |mJy                 |1.40E+09 |   1.8E-03  |+/-0.7E-03|Jy|2007MNRAS.380..199I|rms uncertainty|       1.4 GHz       | Broad-band measurement|10 52 28.995 +57 22 22.42 (J2000)| Flux integrated from map|                                        |From reprocessed raw data
