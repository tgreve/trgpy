
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-04-05T08:15:36PDT



Photometric Data for SMMJ021738-050339a, z=2.037

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|250 microns (SPIRE) | 18.2     |+/-3.6  |mJy |1.199e+12|18.2E-03  |+/-3.6E-03  |Jy|Reference          |uncertainty       | | | | |
2|350 microns (SPIRE) | 17.0     |+/-4.2  |mJy |8.57e+11|17.0E-03   |+/-4.2E-03  |Jy|Reference          |uncertainty       | | | | |
3|500 microns (SPIRE) | 10.9     |+/-4.8  |mJy |5.996e+11|10.9E-03  |+/-4.8E-03  |Jy|Reference          |uncertainty       | | | | |
1|850 microns (SCUBA) | 2.2      |+/-0.85 |mJy   |3.53E+11|2.2E-03|+/-0.85E-03|Jy|2004ApJ...614..671C|1 sigma|       850 microns   | Broad-band measurement|163656.28 +405912.2 (J2000)| Flux integrated from map|                                        |From new raw data
2|2.0 mm (PdBI)       | 0.4      |+/-0.1  |mJy   |1.54E+11|0.4E-03|+/-0.1E-03|Jy|2010Natur.464..733S|uncertainty|       2.8 microns   | Broad-band measurement|21 35 11.6 -01 02 52.0 (J2000)| Flux in fixed aperture|                                        |From new raw data
6|1.4 GHz (VLA)       | 92.5     |+/-12   |uJy |1.40E+09|92.5E-06|+/-12.E-06|Jy|2006MNRAS.371..963B|1 sigma|       1.4 GHz       | Broad-band measurement|16 36 55.767 +40 59 09.97 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
