
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-06-16T05:28:49PDT



Photometric Data for CFRS 14.0711

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|F606W (total)       | 22.79     |+/-0.06 |mag                 |5.05E+14|  2.60E-06|+/-1.48E-07|Jy|2002ApJS..142....1S|68% confidence|5934       A         | Broad-band measurement|141756.838 +523159.62 (J2000)| Flux integrated from map|                                        |From new raw data
2|V (HST/F606W)       | 22.74     ||mag                 |5.05E+14|  2.73E-06||Jy|2005ApJS..159...41V|no uncertainty reported|    5934   A         | Broad-band measurement|14 17 56.832 +52 31 59.60 (J2000)| Flux in fixed aperture|1.5" diameter aperture                  |From new raw data
3|V (HST/F606W)       | 22.37     ||mag                 |5.05E+14|  3.83E-06||Jy|2005ApJS..159...41V|no uncertainty reported|    5934   A         | Broad-band measurement|14 17 56.832 +52 31 59.60 (J2000)| Total flux|Magnitude measured with FOCAS           |From new raw data
4|V (HST/F606W)       | 21.87     ||mag                 |5.05E+14|  6.07E-06||Jy|2005ApJS..159...41V|no uncertainty reported|    5934   A         | Broad-band measurement|14 17 56.832 +52 31 59.60 (J2000)| Total flux|Magnitude measured with GIM2D           |From new raw data
5|F606W (HST)         | 22.30     || mag                |5.05E+14|  4.09E-06||Jy|2004A&A...421..847Z|no uncertainty reported|    5934   A         | Broad-band measurement|| Flux in fixed aperture|3" aperture                             |From reprocessed raw data
6|I (HST/F814W)       | 21.73     ||mag                 |3.78E+14|  5.06E-06||Jy|2005ApJS..159...41V|no uncertainty reported|    7924   A         | Broad-band measurement|14 17 56.832 +52 31 59.60 (J2000)| Flux in fixed aperture|1.5" diameter aperture                  |From new raw data
7|I (HST/F814W)       | 21.33     ||mag                 |3.78E+14|  7.32E-06||Jy|2005ApJS..159...41V|no uncertainty reported|    7924   A         | Broad-band measurement|14 17 56.832 +52 31 59.60 (J2000)| Total flux|Magnitude measured with FOCAS           |From new raw data
8|I (HST/F814W)       | 22.78     ||mag                 |3.78E+14|  1.92E-06||Jy|2005ApJS..159...41V|no uncertainty reported|    7924   A         | Broad-band measurement|14 17 56.832 +52 31 59.60 (J2000)| Total flux|Magnitude measured with GIM2D           |From new raw data
9|F814W (total)       | 21.87     |+/-0.04 |mag                 |3.78E+14|  4.45E-06|+/-1.67E-07|Jy|2002ApJS..142....1S|68% confidence|7924       A         | Broad-band measurement|141756.838 +523159.62 (J2000)| Flux integrated from map|                                        |From new raw data
10|F814W (HST)         | 21.24     || mag                |3.78E+14|  7.95E-06||Jy|2004A&A...421..847Z|no uncertainty reported|    7924   A         | Broad-band measurement|| Flux in fixed aperture|3" aperture                             |From reprocessed raw data
11|CO(3-2) (PdBI)      |           |+/-0.13 |Jy km/s             |3.46E+11||+/-7.08E+04|Jy-Hz|2010Natur.463..781T|1 sigma|   345.998 GHz       | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|                                        |From new raw data
