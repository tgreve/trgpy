
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-07-10T12:49:16PDT



Photometric Data for LEDA 2823818

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|H{beta} (VLT)       | 1.9E-15   |+/-0.1E-15|erg/s/cm^2^         |6.17E+14|  1.90E+08|+/-1.00E+07|Jy-Hz|2008A&A...491..407N|uncertainty|      4861 A         | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|                                        |From new raw data
2|[O III] 4959 (VLT)  | 2.2E-15   |+/-0.1E-15|erg/s/cm^2^         |6.05E+14|  2.20E+08|+/-1.00E+07|Jy-Hz|2008A&A...491..407N|uncertainty|      4959 A         | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|                                        |From new raw data
3|[O III] 5007 (VLT)  | 6.6E-15   |+/-0.4E-15|erg/s/cm^2^         |5.99E+14|  6.60E+08|+/-4.00E+07|Jy-Hz|2008A&A...491..407N|uncertainty|      5007 A         | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|                                        |From new raw data
4|[O I] 6300 (VLT)    | 0.74E-15  |+/-0.07E-15|erg/s/cm^2^         |4.76E+14|  7.40E+07|+/-7.00E+06|Jy-Hz|2008A&A...491..407N|uncertainty|      6300 A         | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|                                        |From new raw data
5|H{alpha}+[NII] (VLT)| 9.75E-15  |+/-0.59E-15|erg/s/cm^2^         |4.56E+14|  9.75E+08|+/-5.90E+07|Jy-Hz|2008A&A...491..407N|uncertainty|      6573 A         | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|Flux of blended line                    |From new raw data
6|[S II] (VLT)        | 2.40E-15  |+/-0.16E-15|erg/s/cm^2^         |4.46E+14|  2.40E+08|+/-1.60E+07|Jy-Hz|2008A&A...491..407N|uncertainty|    6723.5 A         | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|Flux of blended line                    |From new raw data
7|3.6 microns (IRAC)  | 40.4      |+/-4.3  | microJy            |8.44E+13|  4.04E-05|+/-4.30E-06|Jy|2007ApJS..171..353S|uncertainty|   3.550   microns   | Broad-band measurement|04 08 51.5 -24 18 16.39 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
8|4.5 microns (IRAC)  | 43.3      |+/-4.6  | microJy            |6.67E+13|  4.33E-05|+/-4.60E-06|Jy|2007ApJS..171..353S|uncertainty|   4.493   microns   | Broad-band measurement|04 08 51.5 -24 18 16.39 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
9|5.8 microns (IRAC)  ||<51.6      | microJy            |5.23E+13||5.16E-05|Jy|2007ApJS..171..353S|3 sigma|   5.731   microns   | Broad-band measurement|04 08 51.5 -24 18 16.39 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
10|8.0 microns (IRAC)  | 63.5      |+/-14.5 | microJy            |3.81E+13|  6.35E-05|+/-1.45E-05|Jy|2007ApJS..171..353S|uncertainty|   7.872   microns   | Broad-band measurement|04 08 51.5 -24 18 16.39 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
11|16 microns (IRS)    | 242.0     |+/-34.6 | microJy            |1.87E+13|  2.42E-04|+/-3.46E-05|Jy|2007ApJS..171..353S|uncertainty|      16   microns   | Broad-band measurement|04 08 51.5 -24 18 16.39 (J2000)| Flux in fixed aperture|6" diameter aperture                    |From reprocessed raw data
12|24 microns (MIPS)   | 1420.0    |+/-83.7 | microJy            |1.27E+13|  1.42E-03|+/-8.37E-05|Jy|2007ApJS..171..353S|uncertainty|   23.68   microns   | Broad-band measurement|04 08 51.5 -24 18 16.39 (J2000)| Flux in fixed aperture|13" diameter aperture                   |From reprocessed raw data
13|70 microns (MIPS)   | 24700     |+/-2306 | microJy            |4.20E+12|  2.47E-02|+/-2.31E-03|Jy|2007ApJS..171..353S|uncertainty|   71.42   microns   | Broad-band measurement|04 08 51.5 -24 18 16.39 (J2000)| Flux in fixed aperture|35" diameter aperture                   |From reprocessed raw data
14|160 microns (MIPS)  ||<47700     | microJy            |1.92E+12||4.77E-02|Jy|2007ApJS..171..353S|3 sigma|   155.9   microns   | Broad-band measurement|04 08 51.5 -24 18 16.39 (J2000)| Flux in fixed aperture|50" diameter aperture                   |From reprocessed raw data
15|4.85 GHz            | 129       |+/-12   |milliJy             |4.85E+09|  1.29E-01|+/-1.20E-02|Jy|1994ApJS...90..179G|rms noise|4.85       GHz       | Broad-band measurement|040850.9 -241819 (J2000)| Modelled datum|                                        |From new raw data; Corrected for contaminating sources
16|1.4GHz (VLA)              | 625.6     |+/-18.8 |milliJy             |1.40E+09|  6.26E-01|+/-1.88E-02|Jy|1998AJ....115.1693C|uncertainty|    1.40   GHz       | Broad-band measurement|04 08 51.38 -24 18 15.3 (J2000)| Flux integrated from map|                                        |From new raw data
17|408 MHz             | 2.92      |+/-0.10 |Jy                  |4.08E+08|  2.92E+00|+/-1.00E-01|Jy|1981MNRAS.194..693L|rms noise|408        MHz       | Broad-band measurement|040644.2 -242613 (B1950)| Modelled datum|                                        |From new raw data; Corrected for contaminating sources
18|365 MHz (Texas)     | 3.881     |+/-0.071|Jy                  |3.65E+08|  3.88E+00|+/-7.10E-02|Jy|1996AJ....111.1945D|internal error|365        MHz       | Broad-band measurement; obtained by interpolation over frequency|040644.358 -242606.43 (B1950)| Integrated from scans|Model:P;MFlag:+;EFlag:+;LFlag:+.        |From new raw data
19|74 MHz (VLA)        | 16.77     |+/-1.71 | Jy                 |7.38E+07|  1.68E+01|+/-1.71E+00|Jy|2007AJ....134.1245C|rms uncertainty|    73.8   MHz       | Broad-band measurement|04 08 51.55 -24 18 13.6 (J2000)| Flux integrated from map|Corrected for clean bias                |From new raw data
