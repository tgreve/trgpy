
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-07-10T07:32:02PDT



Photometric Data for PC 1643+4631A

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|CCD grism r_4       | 20.06     |+/-0.30 |mag                 |4.50E+14|  2.76E-05|+/-8.79E-06|Jy|1994AJ....107.1245S|rms uncertainty|6659       A         | Broad-band measurement; broad-band flux derived by integration over spectrum|164333.5 +463138 (B1950)| Integrated from scans|                                        |From new raw data
