
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-07-08T06:26:59PDT



Photometric Data for MIPS J123644.0+621450.5

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|U (KPNO) AB         | 25.65     ||mag                 |8.44E+14|  2.00E-07||Jy|2006ApJ...653.1004R|no uncertainty reported|    3550   A         | Broad-band measurement|123644.13 +621450.7 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data; derived from aflux in a different band and a color
2|G (KECK) AB         | 24.78     ||mag                 |6.27E+14|  4.45E-07||Jy|2006ApJ...653.1004R|no uncertainty reported|    4780   A         | Broad-band measurement|123644.13 +621450.7 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data; derived from aflux in a different band and a color
3|R (KECK) AB         | 24.25     ||mag                 |4.39E+14|  7.25E-07||Jy|2006ApJ...653.1004R|no uncertainty reported|    6830   A         | Broad-band measurement|123644.13 +621450.7 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data
4|J (WIRC) AB         | 23.16     ||mag                 |2.40E+14|  1.98E-06||Jy|2006ApJ...653.1004R|no uncertainty reported|   1.250   microns   | Broad-band measurement|123644.13 +621450.7 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data
5|K_s (WIRC) AB       | 22.00     ||mag                 |1.39E+14|  5.75E-06||Jy|2006ApJ...653.1004R|no uncertainty reported|   2.150   microns   | Broad-band measurement|123644.13 +621450.7 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data
6|3.6 microns IRAC AB | 21.42     |+/-0.07 |mag                 |8.44E+13|  9.82E-06|+/-6.33E-07|Jy|2006ApJ...653.1004R|uncertainty|   3.550   microns   | Broad-band measurement|123644.13 +621450.7 (J2000)| Flux integrated from map|                                        |From new raw data
7|4.5 microns IRAC AB | 21.26     |+/-0.07 |mag                 |6.67E+13|  1.14E-05|+/-7.33E-07|Jy|2006ApJ...653.1004R|uncertainty|   4.493   microns   | Broad-band measurement|123644.13 +621450.7 (J2000)| Flux integrated from map|                                        |From new raw data
8|5.8 microns IRAC AB | 21.25     |+/-0.11 |mag                 |5.23E+13|  1.15E-05|+/-1.16E-06|Jy|2006ApJ...653.1004R|uncertainty|   5.731   microns   | Broad-band measurement|123644.13 +621450.7 (J2000)| Flux integrated from map|                                        |From new raw data
9|8.0 microns IRAC AB | 21.62     |+/-0.21 |mag                 |3.81E+13|  8.17E-06|+/-1.58E-06|Jy|2006ApJ...653.1004R|uncertainty|   7.872   microns   | Broad-band measurement|123644.13 +621450.7 (J2000)| Flux integrated from map|                                        |From new raw data
10|24 microns (MIPS)   | 143.9     |+/-4.1  |microJy             |1.27E+13|  1.44E-04|+/-4.10E-06|Jy|2011A&A...528A..35M|uncertainty|     23.68 microns   | Broad-band measurement|12 36 44.03 +62 14 50.48 (J2000)| Flux integrated from map|                                        |From new raw data
1|24 microns (MIPS)   | 123       |+/-29   |microJy             |1.27E+13|123.E-06|29.0E-06|Jy|2009ApJ...694.1517D|3sigma uncertainty|     23.68 microns   | Broad-band measurement|12 37 11.89 +62 22 11.8 (J2000)| Flux integrated from map|                                        |From new raw data
11|70 microns (MIPS)   ||<4.7       |milliJy             |4.20E+12||4.70E-03|Jy|2011A&A...528A..35M|no uncertainty reported|     71.42 microns   | Broad-band measurement|12 36 44.03 +62 14 50.48 (J2000)| Flux integrated from map|                                        |From new raw data
2|70 microns (MIPS)   |           |<2.7    |mJy             |4.20E+12|        |2.7E-03|Jy|2009ApJ...699.1610H|3 sigma|     71.42 microns   | Broad-band measurement|221804.42 +002154.4 (J2000)| Flux in fixed aperture|                                        |From new raw data
12|340 GHz (SMA)       | 5.27      |+/-1.14 |milliJy             |3.40E+11|  5.27E-03|+/-1.14E-03|Jy|2011ApJ...726L..18W|uncertainty|       340 GHz       | Broad-band measurement|189.18324 62.24741 (J2000)| Flux integrated from map|Primary beam corrected                  |From new raw data
3|850 microns (SCUBA) |           |<9.4    |mJy             |3.53E+11|        |9.4E-03|Jy|2005MNRAS.358..149P|3sigma uncertainty|     850   microns   | Broad-band measurement|12 37 11.7 +62 22 12 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
4|1200 microns (MAMBO)|           |<4.2    |mJy             |2.50E+11|        |4.2E-03|Jy|2004MNRAS.354..779G|3sigma uncertainty|      1200 microns   | Broad-band measurement|16 36 55.9 +40 59 12 (J2000)| Flux integrated from map|S/N = 3.66                              |From new raw data
13|1.4 GHz (VLA)       | 32.6      |+/-7.3  |microJy             |1.40E+09|  3.26E-05|+/-7.30E-06|Jy|2010ApJS..188..178M|uncertainty|       1.4 GHz       | Broad-band measurement|12 36 44.01 +62 14 50.5 (J2000)| Total flux; Beam filling or dilution corrected|Major=0.5"; Minor=0.0"; PA=135 deg      |From new raw data
5|1.4 GHz (VLA)       | 39.6      |+/-8.7  | microJy        |1.40E+09| 39.6E-06|+/-8.7E-06|Jy|2006MNRAS.371..963B|1 sigma|       1.4 GHz       | Broad-band measurement|16 36 55.767 +40 59 09.97 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
