
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-06-11T07:56:28PDT



Photometric Data for BzK16000 (z=1.522)

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|R (Keck II) AB      | 23.61     | | mag                |4.62E+14|  1.31E-06| |Jy|2004AJ....127.3121W|no uncertainty reported|   648.7   A         | Broad-band measurement|12 36 30.079 +62 14 28.03 (J2000)| Total flux|                                        |From new raw data
2|H{alpha} (Subaru)   | 17.4E-17  |+/-4.8E-17|erg/s/cm^2^         |4.57E+14|  1.74E+07|+/-4.80E+06|Jy-Hz|2010ApJ...718..112Y|uncertainty|      6563 A         | Line measurement; flux integrated over line; lines measured in emission|12 36 30.08 +62 14 27.9 (J2000)| Flux integrated from map|                                        |From new raw data
3|K_s (Subaru) AB     | 20.6      | |mag                 |1.39E+14|  2.09E-05| |Jy|2010ApJ...718..112Y|no uncertainty reported|      2.15 microns   | Broad-band measurement|12 36 30.08 +62 14 27.9 (J2000)| Total flux|                                        |Averaged from previously published data
4|3.6 microns (IRAC)  | 41.00     |+/-2.05 |microJy             |8.44E+13|  4.10E-05|+/-2.05E-06|Jy|2011AJ....141....1T|rms uncertainty|     3.550 microns   | Broad-band measurement|189.125366 62.241077 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
5|4.5 microns (IRAC)  | 43.40     |+/-2.17 |microJy             |6.67E+13|  4.34E-05|+/-2.17E-06|Jy|2011AJ....141....1T|rms uncertainty|     4.493 microns   | Broad-band measurement|189.125366 62.241077 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
6|5.8 microns (IRAC)  | 34.20     |+/-1.75 |microJy             |5.23E+13|  3.42E-05|+/-1.75E-06|Jy|2011AJ....141....1T|rms uncertainty|     5.731 microns   | Broad-band measurement|189.125366 62.241077 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
7|8.0 microns (IRAC)  | 29.00     |+/-1.52 |microJy             |3.81E+13|  2.90E-05|+/-1.52E-06|Jy|2011AJ....141....1T|rms uncertainty|     7.872 microns   | Broad-band measurement|189.125366 62.241077 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
8|16 microns (IRS)    | 111.0     |+/-8.7  |microJy             |1.90E+13|  1.11E-04|+/-8.70E-06|Jy|2011AJ....141....1T|rms uncertainty|      15.8 microns   | Broad-band measurement|189.125366 62.241077 (J2000)| From fitting to map|                                        |From new raw data
9|24 microns (MIPS)   | 188.0     |+/-5.8  |microJy             |1.27E+13|  1.88E-04|+/-5.80E-06|Jy|2011AJ....141....1T|rms uncertainty|     23.68 microns   | Broad-band measurement|189.125366 62.241077 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
10|24 microns (MIPS)  | 190.0     |+/-6.0  |microJy             |1.27E+13|  1.90E-04|+/-6.0E-06|Jy|2011AJ....141....1T|rms uncertainty|     23.68 microns   | Broad-band measurement|189.125366 62.241077 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
11|70 microns (PACS)  |           |<2.0    |mJy                 |4.283E+12|         |2.0E-03|Jy|2004MNRAS.354..779G|3sigma uncertainty|      1200 microns   | Broad-band measurement|16 36 55.9 +40 59 12 (J2000)| Flux integrated from map|S/N = 3.66                              |From new raw data
12|100 microns (PACS) | 1.6       |+/-0.6  |microJy             |2.998e+12| 1.6E-03 |+/-0.6E-03 |Jy|2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
13|160 microns (PACS) | 3.7       |+/-0.9  |microJy             |1.874e+12| 3.7E-03 |+/-0.9E-03 |Jy|2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
14|250 microns (SPIRE)| 9.2       |+/-2.5  |mJy                 |1.199e+12| 9.2E-03 |+/-2.5e-03 |Jy|2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
15|350 microns (SPIRE)|           |<9.0    |mJy                 |8.565E+11|         |9.0E-03|Jy|2004MNRAS.354..779G|3sigma uncertainty|      1200 microns   | Broad-band measurement|16 36 55.9 +40 59 12 (J2000)| Flux integrated from map|S/N = 3.66                              |From new raw data
16|500 microns (SPIRE)|           |<12.0   |mJy                 |5.996E+11|         |12.0E-03|Jy|2004MNRAS.354..779G|3sigma uncertainty|      1200 microns   | Broad-band measurement|16 36 55.9 +40 59 12 (J2000)| Flux integrated from map|S/N = 3.66                              |From new raw data
17|1160 microns (Penner)|         |<1.7    |mJy                 |2.58442E+11|       |1.7E-03|Jy|2004MNRAS.354..779G|3sigma uncertainty|      1200 microns   | Broad-band measurement|16 36 55.9 +40 59 12 (J2000)| Flux integrated from map|S/N = 3.66                              |From new raw data
18|45.6 GHz (VLA)     |           |<360.   |microJy             |45.6E+09|          |360.E-06|Jy|2006MNRAS.371..963B|2sigma|       1.4 GHz       | Broad-band measurement|16 36 55.767 +40 59 09.97 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
19|1.4 GHz (VLA)      | 19.0      |+/-6.0  |microJy             |1.40E+09| 19.0E-06|+/-6.0E-06|Jy|2006MNRAS.371..963B|1 sigma|       1.4 GHz       | Broad-band measurement|16 36 55.767 +40 59 09.97 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
