
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-05-28T01:50:15PDT



Photometric Data for PJ160917.8, z=3.2553

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
2|J (2MASS)           | 0.05     |+/-0.15 |mag          |2.40E+14|  0.05E-03|+/-0.15E-03|Jy|2004ApJ...616...71S|1 sigma|    1.25   microns   | Broad-band measurement| | Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
1|H_total (2MASS)     | 0.89    |+/-0.09|mag            |1.82E+14|  0.89E-03|+/-0.09E-04|Jy|20032MASX.C.......:|1 sigma uncert.| 1.65      microns   | Broad-band measurement|041437.75 +053442.6 (J2000)| Total flux|                                        |From new raw data
3|K_s_ (2MASS)        | 0.68     |+/-0.11 |mag          |1.38E+14|  0.68E-03|+/-0.11E-03|Jy|2004ApJ...616...71S|1 sigma|    2.17   microns   | Broad-band measurement| | Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
26|22 microns (WISE)  |        |<5.4|mJy            |1.36E+13||5.4E-03|Jy|2012AJ....144...49W|3sigma limit|        22 microns   | Broad-band measurement|213.942657 +11.495400 (J2000)| Not reported in paper|                                        |Averaged from previously published data
1|250 microns (SPIRE) | 568.0     |+/-57.  |mJy         |1.199e+12|568.0E-03 |+/-57.0e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
1|250 microns (SPIRE) | 765.0     |+/-7.  |mJy         |1.199e+12|765.0E-03 |+/-7.0e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
3|350 microns (SPIRE) | 693.0     |+/-69.  |mJy         |8.565e+11|693.0E-03 |+/-69.0e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
3|350 microns (SPIRE) | 865.0     |+/-8.  |mJy         |8.565e+11|865.0E-03 |+/-8.0e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
5|350 microns (PLANCK) | 1083.0    |+/-255.  |mJy       |8.57e+11|1083.0E-03 |+/-255.0e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
5|500 microns (SPIRE) | 512.0     |+/-51.  |mJy         |5.996e+11|512.0E-03 |+/-51.0e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
5|500 microns (SPIRE) | 696.0     |+/-7.  |mJy         |5.996e+11|696.0E-03 |+/-7.0e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
9|850 microns (SCUBA) | 191.0     |+/-16. |milliJy       |3.53E+11|  191.E-03|+/-16.E-03 |Jy|2002MNRAS.331..495S|no uncertainty reported|     850   microns   | Broad-band measurement|140105.0 +025225 (J2000)| Flux integrated from map|                                        |From new raw data
2|1.1mm (AzTEC)        | 73.8     |+/-7.0  | mJy        |2.73E11| 73.8E-3| 7.0E-3 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
5|GISMO(2000.0um)     |  8.4   |+/-0.6 |mJy          |150.000E+9|8.4E-03 |+/-0.6E-03|Jy|2010ApJ...709..210K|uncertainty|      870  microns   | Broad-band measurement|16 35 55.67 +66 12 59.51 (J2000)| Flux integrated from map|                                        |From new raw data
5|VLA Ka-band 31.1GHz|  230   |+/-20 |mJy          |31.056E+9|230.0E-06 |+/-20E-06|Jy|2010ApJ...709..210K|uncertainty|      870  microns   | Broad-band measurement|16 35 55.67 +66 12 59.51 (J2000)| Flux integrated from map|                                        |From new raw data
5|VLA K-band 23.2GHz    |  303   |+/-14 |mJy          |23.1991E+9|303.0E-06 |+/-14E-06|Jy|2010ApJ...709..210K|uncertainty|      870  microns   | Broad-band measurement|16 35 55.67 +66 12 59.51 (J2000)| Flux integrated from map|                                        |From new raw data
21|1.4GHz (VLA)       |   1.5 |+/-0.3|mJy| 1.4E9   |1.5E-03 |0.3E-03 |Jy |2003MNRAS.343..293M|3rms uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
