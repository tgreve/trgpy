
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-06-16T05:23:52PDT



Photometric Data for SDSS J141642.10+522519.2

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|u (SDSS PSF) AB     | 23.215    |+/-0.671|asinh mag           |8.36E+14|  1.81E-06|+/-1.29E-06|Jy|2007SDSS6.C...0000:|based on count statistics only|3585       A         | Broad-band measurement|214.1754254556 52.4220134483 (J2000)| Modelled datum|SDSS flags: CANONICAL_CENTER - used canonical, not local, center; NOPETRO - no Petrosian radius could be determined; NOPETRO_BIG - Petrosian radius is larger than extracted radial profile; MANYR50 - more than one 50% radius; BAD_RADIAL - some low S/N radial points; ELLIPFAINT - no isophotal fits performed; AMOMENT_FAINT - too faint for adaptive moments;|From new raw data
2|u (SDSS CModel) AB  | 22.889    ||asinh mag           |8.36E+14|  2.53E-06||Jy|2007SDSS6.C...0000:|no uncertainty reported|3585       A         | Broad-band measurement|214.1754254556 52.4220134483 (J2000)| Modelled datum|SDSS flags: CANONICAL_CENTER - used canonical, not local, center; NOPETRO - no Petrosian radius could be determined; NOPETRO_BIG - Petrosian radius is larger than extracted radial profile; MANYR50 - more than one 50% radius; BAD_RADIAL - some low S/N radial points; ELLIPFAINT - no isophotal fits performed; AMOMENT_FAINT - too faint for adaptive moments;|From new raw data
3|u (SDSS Model) AB   | 23.148    |+/-0.853|asinh mag           |8.36E+14|  1.94E-06|+/-1.73E-06|Jy|2007SDSS6.C...0000:|based on count statistics only|3585       A         | Broad-band measurement|214.1754254556 52.4220134483 (J2000)| Modelled datum|SDSS flags: CANONICAL_CENTER - used canonical, not local, center; NOPETRO - no Petrosian radius could be determined; NOPETRO_BIG - Petrosian radius is larger than extracted radial profile; MANYR50 - more than one 50% radius; BAD_RADIAL - some low S/N radial points; ELLIPFAINT - no isophotal fits performed; AMOMENT_FAINT - too faint for adaptive moments;|From new raw data
4|g (SDSS PSF) AB     | 23.350    |+/-0.250|asinh mag           |6.17E+14|  1.60E-06|+/-3.97E-07|Jy|2007SDSS6.C...0000:|based on count statistics only|4858       A         | Broad-band measurement|214.1754254556 52.4220134483 (J2000)| Modelled datum|SDSS flags: CANONICAL_CENTER - used canonical, not local, center; NOPETRO - no Petrosian radius could be determined; BAD_RADIAL - some low S/N radial points; PETROFAINT - Petrosian radius measured at very low surface brightness; ELLIPFAINT - no isophotal fits performed; AMOMENT_FAINT - too faint for adaptive moments;|From new raw data
5|g (SDSS CModel) AB  | 22.179    ||asinh mag           |6.17E+14|  4.86E-06||Jy|2007SDSS6.C...0000:|no uncertainty reported|4858       A         | Broad-band measurement|214.1754254556 52.4220134483 (J2000)| Modelled datum|SDSS flags: CANONICAL_CENTER - used canonical, not local, center; NOPETRO - no Petrosian radius could be determined; BAD_RADIAL - some low S/N radial points; PETROFAINT - Petrosian radius measured at very low surface brightness; ELLIPFAINT - no isophotal fits performed; AMOMENT_FAINT - too faint for adaptive moments;|From new raw data
6|g (SDSS Model) AB   | 22.842    |+/-0.216|asinh mag           |6.17E+14|  2.61E-06|+/-5.35E-07|Jy|2007SDSS6.C...0000:|based on count statistics only|4858       A         | Broad-band measurement|214.1754254556 52.4220134483 (J2000)| Modelled datum|SDSS flags: CANONICAL_CENTER - used canonical, not local, center; NOPETRO - no Petrosian radius could be determined; BAD_RADIAL - some low S/N radial points; PETROFAINT - Petrosian radius measured at very low surface brightness; ELLIPFAINT - no isophotal fits performed; AMOMENT_FAINT - too faint for adaptive moments;|From new raw data
7|r (SDSS CModel) AB  | 22.110    ||asinh mag           |4.77E+14|  5.16E-06||Jy|2007SDSS6.C...0000:|no uncertainty reported|6290       A         | Broad-band measurement|214.1754254556 52.4220134483 (J2000)| Modelled datum|SDSS flags: NOPETRO - no Petrosian radius could be determined; MANYR90 - more than one 90% radius; BAD_RADIAL - some low S/N radial points; PETROFAINT - Petrosian radius measured at very low surface brightness; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding; CANONICAL_BAND - this band was primary (usually r);|From new raw data
8|r (SDSS PSF) AB     | 22.507    |+/-0.172|asinh mag           |4.77E+14|  3.56E-06|+/-5.80E-07|Jy|2007SDSS6.C...0000:|based on count statistics only|6290       A         | Broad-band measurement|214.1754254556 52.4220134483 (J2000)| Modelled datum|SDSS flags: NOPETRO - no Petrosian radius could be determined; MANYR90 - more than one 90% radius; BAD_RADIAL - some low S/N radial points; PETROFAINT - Petrosian radius measured at very low surface brightness; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding; CANONICAL_BAND - this band was primary (usually r);|From new raw data
9|r (SDSS Model) AB   | 22.110    |+/-0.168|asinh mag           |4.77E+14|  5.16E-06|+/-8.10E-07|Jy|2007SDSS6.C...0000:|based on count statistics only|6290       A         | Broad-band measurement|214.1754254556 52.4220134483 (J2000)| Modelled datum|SDSS flags: NOPETRO - no Petrosian radius could be determined; MANYR90 - more than one 90% radius; BAD_RADIAL - some low S/N radial points; PETROFAINT - Petrosian radius measured at very low surface brightness; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding; CANONICAL_BAND - this band was primary (usually r);|From new raw data
10|i (SDSS PSF) AB     | 22.058    |+/-0.164|asinh mag           |3.89E+14|  5.38E-06|+/-8.36E-07|Jy|2007SDSS6.C...0000:|based on count statistics only|7706       A         | Broad-band measurement|214.1754254556 52.4220134483 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; ELLIPFAINT - no isophotal fits performed; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
11|i (SDSS CModel) AB  | 21.657    ||asinh mag           |3.89E+14|  7.84E-06||Jy|2007SDSS6.C...0000:|no uncertainty reported|7706       A         | Broad-band measurement|214.1754254556 52.4220134483 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; ELLIPFAINT - no isophotal fits performed; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
12|i (SDSS Model) AB   | 21.736    |+/-0.179|asinh mag           |3.89E+14|  7.28E-06|+/-1.22E-06|Jy|2007SDSS6.C...0000:|based on count statistics only|7706       A         | Broad-band measurement|214.1754254556 52.4220134483 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; ELLIPFAINT - no isophotal fits performed; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
13|z (SDSS PSF) AB     | 21.179    |+/-0.245|asinh mag           |3.25E+14|  1.15E-05|+/-2.85E-06|Jy|2007SDSS6.C...0000:|based on count statistics only|9222       A         | Broad-band measurement|214.1754254556 52.4220134483 (J2000)| Modelled datum|SDSS flags: CANONICAL_CENTER - used canonical, not local, center; MANYR50 - more than one 50% radius; MANYR90 - more than one 90% radius; BAD_RADIAL - some low S/N radial points; INTERP - object contains interpolated-over pixels; ELLIPFAINT - no isophotal fits performed;|From new raw data
14|z (SDSS CModel) AB  | 20.031    ||asinh mag           |3.25E+14|  3.44E-05||Jy|2007SDSS6.C...0000:|no uncertainty reported|9222       A         | Broad-band measurement|214.1754254556 52.4220134483 (J2000)| Modelled datum|SDSS flags: CANONICAL_CENTER - used canonical, not local, center; MANYR50 - more than one 50% radius; MANYR90 - more than one 90% radius; BAD_RADIAL - some low S/N radial points; INTERP - object contains interpolated-over pixels; ELLIPFAINT - no isophotal fits performed;|From new raw data
15|z (SDSS Model) AB   | 20.987    |+/-0.307|asinh mag           |3.25E+14|  1.39E-05|+/-4.20E-06|Jy|2007SDSS6.C...0000:|based on count statistics only|9222       A         | Broad-band measurement|214.1754254556 52.4220134483 (J2000)| Modelled datum|SDSS flags: CANONICAL_CENTER - used canonical, not local, center; MANYR50 - more than one 50% radius; MANYR90 - more than one 90% radius; BAD_RADIAL - some low S/N radial points; INTERP - object contains interpolated-over pixels; ELLIPFAINT - no isophotal fits performed;|From new raw data
16|K_s (Keck)          | 17.74     || mag                |1.39E+14|  4.97E-05||Jy|2007MNRAS.382..109T|no uncertainty reported|      2.15 microns   | Broad-band measurement|214.17549 +52.42204 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
