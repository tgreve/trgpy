

Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.


queryDateTime:2009-11-03T15:07:35PST






Photometric Data for MIPS506 (z=2.4704)

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
4|R (KPNO)            | 1.237     ||microJy             |4.66E+14|  1.24E-06||Jy|2007ApJ...658..778Y|no uncertainty reported|    6440   A         | Broad-band measurement|171138.59 +583836.7 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data
5|R (Cousins) m_aper  | 23.41     |+/-0.06 |mag                 |4.65E+14|  1.32E-06|+/-7.31E-08|Jy|2004AJ....128....1F|based on count statistics only|6440       A         | Broad-band measurement|171138.688 +583836.38 (J2000)| Flux in fixed aperture|3-arcsecond aperture                    |From new raw data
6|R (Cousins) m_tot   | 23.44     |+/-0.08 |mag                 |4.65E+14|  1.29E-06|+/-9.49E-08|Jy|2004AJ....128....1F|based on count statistics only|6440       A         | Broad-band measurement|171138.688 +583836.38 (J2000)| Total flux|                                        |From new raw data
7|F160W (HST NICMOS)  | 20.78     ||mag                 |1.87E+14|  5.09E-06||Jy|2011ApJ...730..125Z|no uncertainty reported|      1.60 microns   | Broad-band measurement|| Flux integrated from map|                                        |From new raw data
8|F160W (HST NICMOS)  | 21.66     || mag                |1.86E+14|  2.26E-06||Jy|2008ApJ...680..232D|no uncertainty reported|      1.61 microns   | Broad-band measurement|17 11 38.52 +58 38 38.58 (J2000)| Flux integrated from map|                                        |From new raw data
9|3.6 microns (IRAC)  | 18        |+/-3    | microJy            |8.44E+13|  1.80E-05|+/-3.00E-06|Jy|2007ApJ...664..713S|uncertainty|   3.550   microns   | Broad-band measurement|| Flux in fixed aperture|7.3" diameter aperture                  |From reprocessed raw data
10|4.5 microns (IRAC)  | 16        |+/-1    | microJy            |6.67E+13|  1.60E-05|+/-1.00E-06|Jy|2007ApJ...664..713S|uncertainty|   4.493   microns   | Broad-band measurement|| Flux in fixed aperture|7.3" diameter aperture                  |From reprocessed raw data
11|5.8 microns (IRAC)  | 26        |+/-18   | microJy            |5.23E+13|  2.60E-05|+/-1.80E-05|Jy|2007ApJ...664..713S|uncertainty|   5.731   microns   | Broad-band measurement|| Flux in fixed aperture|7.3" diameter aperture                  |From reprocessed raw data
14|8.0 microns (IRAC)  | 13        |+/-19   | microJy            |3.81E+13|  1.30E-05|+/-1.90E-05|Jy|2007ApJ...664..713S|uncertainty|   7.872   microns   | Broad-band measurement|| Flux in fixed aperture|7.3" diameter aperture                  |From reprocessed raw data
15|8.0 microns (IRAC)  | 20.000    ||microJy             |3.81E+13|  2.00E-05||Jy|2007ApJ...658..778Y|no uncertainty reported|   7.872   microns   | Broad-band measurement|171138.59 +583836.7 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data
1|MIPS 24um           | 1.06     |+/-0.32 |milliJy             |1.27E+13|  1.06E-03|+/-0.32E-03 |Jy|1996AJ....111.1431B|uncertainty|1.49       GHz       | Broad-band measurement| | Peak flux|                                        |From new raw data
17|24 microns (MIPS)   | 920.141   ||microJy             |1.27E+13|  9.20E-04||Jy|2007ApJ...658..778Y|no uncertainty reported|   23.68   microns   | Broad-band measurement|171138.59 +583836.7 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data; measurementmodified from published value
2|MIPS 70um           |          |<4.5    |milliJy             |4.20E+12|          |4.5E-03|Jy|2010Natur.464..733S|3sigma uncertainty|     71.42 microns   | Broad-band measurement|21 35 11.6 -01 02 52.0 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
18|70 microns (MIPS)   | 7.5       |+/-1.2  | milliJy            |4.20E+12|  7.50E-03|+/-1.20E-03|Jy|2007ApJ...664..713S|estimated error|   71.42   microns   | Broad-band measurement|| Flux in fixed aperture|3 pixel radius aperture                 |From reprocessed raw data
3|MIPS 160um          |          |<30     |milliJy             |1.92E+12|          |30.0E-03|Jy|2009A&A...502..541E|3 sigma|     155.9 microns   | Broad-band measurement| | Flux in fixed aperture|                                        |From reprocessed raw data
4|MAMBO 1200um        | 1.37     |+/-0.53 |milliJy             |2.50E+11|  1.37E-03|+/-0.53E-03|Jy|2004MNRAS.354..779G|3sigma uncertainty|      1200 microns   | Broad-band measurement|16 37 06.7 +40 53 15 (J2000)| Flux integrated from map|S/N = 3.81                              |From new raw data
5|VLA 1.4GHz          | 0.14     |+/-0.03 |milliJy             |1.4E9   |  0.14E-3|+/-0.03E-3|Jy |2003MNRAS.343..293M|3sigma uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
