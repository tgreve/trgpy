
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-07-10T09:29:26PDT



Photometric Data for LEDA 2823016

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|12 microns (ISOCAM) | 1.8       |+/-0.3  |milliJy             |2.50E+13|  1.80E-03|+/-3.00E-04|Jy|2004A&A...421..129S|1 sigma|    12.0   microns   | Broad-band measurement|| From multi-aperture data|                                        |From reprocessed raw data; OBJ_NAME modified from publishedvalue
2|4.85 GHz            | 66        |+/-11   |milliJy             |4.85E+09|  6.60E-02|+/-1.10E-02|Jy|1994ApJS...90..179G|rms noise|4.85       GHz       | Broad-band measurement|021418.7 -115810 (J2000)| Modelled datum|                                        |From new raw data; Corrected for contaminating sources
3|1.4GHz              | 230.4     |+/-8.1  |milliJy             |1.40E+09|  2.30E-01|+/-8.10E-03|Jy|1998AJ....115.1693C|uncertainty|    1.40   GHz       | Broad-band measurement|02 14 17.44 -11 58 45.7 (J2000)| Flux integrated from map|                                        |From new raw data
4|408 MHz             | 1.02      |+/-0.04 |Jy                  |4.08E+08|  1.02E+00|+/-4.00E-02|Jy|1981MNRAS.194..693L|rms noise|408        MHz       | Broad-band measurement|021151.6 -121252 (B1950)| Modelled datum|                                        |From new raw data; Corrected for contaminating sources
5|365 MHz (Texas)     | 1.012     |+/-0.031|Jy                  |3.65E+08|  1.01E+00|+/-3.10E-02|Jy|1996AJ....111.1945D|internal error|365        MHz       | Broad-band measurement; obtained by interpolation over frequency|021151.471 -121243.46 (B1950)| Integrated from scans|Model:P;MFlag:+;EFlag:+;LFlag:+.        |From new raw data
6|74 MHz (VLA)        | 5.03      |+/-0.54 | Jy                 |7.38E+07|  5.03E+00|+/-5.40E-01|Jy|2007AJ....134.1245C|rms uncertainty|    73.8   MHz       | Broad-band measurement|02 14 17.59 -11 58 47.7 (J2000)| Flux integrated from map|Corrected for clean bias                |From new raw data
