
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-07-10T06:33:32PDT



Photometric Data for SDSS J121804.56+470850.1

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|0.5-2 keV           | 2.36E-14  |+/-1.15E-14|erg cm^-2^ s^-1^    |3.02E+17|  7.81E-09|+/-3.81E-09|Jy|2005MNRAS.360..610S|uncertainty|    1.25   keV       | Broad-band measurement|12 18 04.54 +47 08 51.0 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data;Extinction-corrected for Milky Way; NED frequency assigned tomid-point of band in keV
2|FUV (GALEX) AB      ||>23.1173   |mag                 |1.95E+15||2.06E-06|Jy|2012GMSC..C...0000S|3 sigma|1538.6     A         | Broad-band measurement|184.51885663295 47.147693241402 (J2000)| Flux integrated from map|upper limit inside NUV Kron aperture    |From new raw data
3|FUV (GALEX) AB      | 25.3757   |+/-0.944741|mag                 |1.95E+15|  2.57E-07|+/-2.23E-07|Jy|2012GMSC..C...0000S|uncertainty|1538.6     A         | Broad-band measurement|184.51885663295 47.147693241402 (J2000)| Flux in fixed aperture|Flux in 7.5 arcsec diameter aperture    |From new raw data
4|NUV (GALEX) AB      | 22.7827   |+/-0.189429|mag                 |1.29E+15|  2.80E-06|+/-4.88E-07|Jy|2012GMSC..C...0000S|uncertainty|2315.7     A         | Broad-band measurement|184.51885663295 47.147693241402 (J2000)| Flux integrated from map|Kron flux in elliptical aperture        |From new raw data
5|NUV (GALEX) AB      | 23.4039   |+/-0.153309|mag                 |1.29E+15|  1.58E-06|+/-2.23E-07|Jy|2012GMSC..C...0000S|uncertainty|2315.7     A         | Broad-band measurement|184.51885663295 47.147693241402 (J2000)| Flux in fixed aperture|Flux in 7.5 arcsec diameter aperture    |From new raw data
6|u (SDSS PSF) AB     | 21.148    |+/-0.095|asinh mag           |8.36E+14|  1.31E-05|+/-1.15E-06|Jy|2007SDSS6.C...0000:|based on count statistics only|3585       A         | Broad-band measurement|184.5190021705 47.1472503580 (J2000)| Modelled datum|SDSS flags: CHILD - object is part of a blended parent object; BAD_RADIAL - some low S/N radial points; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding; BRIGHTEST_GALAXY_CHILD - brightest child among one parent's children;|From new raw data
7|g (SDSS PSF) AB     | 20.321    |+/-0.023|asinh mag           |6.17E+14|  2.70E-05|+/-5.72E-07|Jy|2007SDSS6.C...0000:|based on count statistics only|4858       A         | Broad-band measurement|184.5190021705 47.1472503580 (J2000)| Modelled datum|SDSS flags: CHILD - object is part of a blended parent object; BAD_RADIAL - some low S/N radial points; BINNED1 - detected at >=5 sigma in original imaging frame;|From new raw data
8|r (SDSS PSF) AB     | 20.034    |+/-0.025|asinh mag           |4.77E+14|  3.52E-05|+/-8.10E-07|Jy|2007SDSS6.C...0000:|based on count statistics only|6290       A         | Broad-band measurement|184.5190021705 47.1472503580 (J2000)| Modelled datum|SDSS flags: CHILD - object is part of a blended parent object; BAD_RADIAL - some low S/N radial points; BINNED1 - detected at >=5 sigma in original imaging frame; CANONICAL_BAND - this band was primary (usually r);|From new raw data
9|i (SDSS PSF) AB     | 19.951    |+/-0.041|asinh mag           |3.89E+14|  3.80E-05|+/-1.43E-06|Jy|2007SDSS6.C...0000:|based on count statistics only|7706       A         | Broad-band measurement|184.5190021705 47.1472503580 (J2000)| Modelled datum|SDSS flags: CHILD - object is part of a blended parent object; BAD_RADIAL - some low S/N radial points; BINNED1 - detected at >=5 sigma in original imaging frame; MAYBE_CR - object may be a cosmic ray;|From new raw data
10|z (SDSS PSF) AB     | 19.786    |+/-0.091|asinh mag           |3.25E+14|  4.33E-05|+/-3.65E-06|Jy|2007SDSS6.C...0000:|based on count statistics only|9222       A         | Broad-band measurement|184.5190021705 47.1472503580 (J2000)| Modelled datum|SDSS flags: CHILD - object is part of a blended parent object; BAD_RADIAL - some low S/N radial points; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding; BRIGHTEST_GALAXY_CHILD - brightest child among one parent's children;|From new raw data
11|450 microns (SCUBA) | 24        |+/-9    |milliJy             |6.66E+11|  2.40E-02|+/-9.00E-03|Jy|2005MNRAS.360..610S|uncertainty|     450   microns   | Broad-band measurement|12 18 04.54 +47 08 51.0 (J2000)| Flux integrated from map|                                        |From new raw data
12|850 microns (SCUBA) | 6.8       |+/-1.2  |milliJy             |3.53E+11|  6.80E-03|+/-1.20E-03|Jy|2005MNRAS.360..610S|uncertainty|     850   microns   | Broad-band measurement|12 18 04.54 +47 08 51.0 (J2000)| Flux integrated from map|Original refcode=2001Sci...294.2516P    |Averaged from previously published data
