

Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.


queryDateTime:2009-11-03T15:07:35PST






Photometric Data for MIPS16080 (z=2.007)

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
4|R (KPNO)            | 2.111     ||microJy             |4.66E+14|  2.11E-06||Jy|2007ApJ...658..778Y|no uncertainty reported|    6440   A         | Broad-band measurement|171844.77 +600115.9 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data
5|R (Cousins) m_tot   | 22.86     |+/-0.05 |mag                 |4.65E+14|  2.20E-06|+/-1.01E-07|Jy|2004AJ....128....1F|based on count statistics only|6440       A         | Broad-band measurement|171844.832 +600116.03 (J2000)| Total flux|                                        |From new raw data
6|R (Cousins) m_aper  | 23.05     |+/-0.04 |mag                 |4.65E+14|  1.84E-06|+/-6.79E-08|Jy|2004AJ....128....1F|based on count statistics only|6440       A         | Broad-band measurement|171844.832 +600116.03 (J2000)| Flux in fixed aperture|3-arcsecond aperture                    |From new raw data
7|F160W (HST NICMOS)         | 20.21     ||mag                 |1.87E+14|  8.60E-06||Jy|2011ApJ...730..125Z|no uncertainty reported|      1.60 microns   | Broad-band measurement|| Flux integrated from map|                                        |From new raw data
8|F160W (HST NICMOS)         | 20.31     || mag                |1.86E+14|  7.84E-06||Jy|2008ApJ...680..232D|no uncertainty reported|      1.61 microns   | Broad-band measurement|17 18 44.83 +60 01 15.82 (J2000)| Flux integrated from map|                                        |From new raw data
10|3.6 microns (IRAC)  | 27        |+/-3    | microJy            |8.44E+13|  2.70E-05|+/-3.00E-06|Jy|2007ApJ...664..713S|uncertainty|   3.550   microns   | Broad-band measurement|| Flux in fixed aperture|7.3" diameter aperture                  |From reprocessed raw data
11|3.6 microns (IRAC)  | 29.98     |+/-4.05 |microJy             |8.42E+13|  3.00E-05|+/-4.05E-06|Jy|2005ApJS..161...41L|uncertainty|3.56       microns   | Broad-band measurement|171844.83 +600115.8 (J2000)| Flux in fixed aperture|Aperture =       4.92 arcsec.           |From new raw data
12|4.5 microns (IRAC)  | 31        |+/-7    | microJy            |6.67E+13|  3.10E-05|+/-7.00E-06|Jy|2007ApJ...664..713S|uncertainty|   4.493   microns   | Broad-band measurement|| Flux in fixed aperture|7.3" diameter aperture                  |From reprocessed raw data
13|4.5 microns (IRAC)  | 31.89     |+/-5.14 |microJy             |6.63E+13|  3.19E-05|+/-5.14E-06|Jy|2005ApJS..161...41L|uncertainty|4.52       microns   | Broad-band measurement|171844.83 +600115.8 (J2000)| Flux in fixed aperture|Aperture =       4.92 arcsec.           |From new raw data
14|5.8 microns (IRAC)  | 38        |+/-24   | microJy            |5.23E+13|  3.80E-05|+/-2.40E-05|Jy|2007ApJ...664..713S|uncertainty|   5.731   microns   | Broad-band measurement|| Flux in fixed aperture|7.3" diameter aperture                  |From reprocessed raw data
15|5.8 microns (IRAC)  ||<100.00    |microJy             |5.23E+13||1.00E-04|Jy|2005ApJS..161...41L|3sigma plate limit|5.73       microns   | Broad-band measurement|171844.83 +600115.8 (J2000)| Flux in fixed aperture|Aperture =       4.92 arcsec.           |From new raw data
18|8.0 microns (IRAC)  | 71        |+/-24   | microJy            |3.81E+13|  7.10E-05|+/-2.40E-05|Jy|2007ApJ...664..713S|uncertainty|   7.872   microns   | Broad-band measurement|| Flux in fixed aperture|7.3" diameter aperture                  |From reprocessed raw data
19|8.0 microns (IRAC)  | 64.978    ||microJy             |3.81E+13|  6.50E-05||Jy|2007ApJ...658..778Y|no uncertainty reported|   7.872   microns   | Broad-band measurement|171844.77 +600115.9 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data
20|8.0 microns (IRAC)  ||<100.00    |microJy             |3.79E+13||1.00E-04|Jy|2005ApJS..161...41L|3sigma plate limit|7.91       microns   | Broad-band measurement|171844.83 +600115.8 (J2000)| Flux in fixed aperture|Aperture =       4.92 arcsec.           |From new raw data
21|8 microns (IRAC) | 1.5       |+/-1   %|milliJy             |3.75E+13|  1.50E-03|+/-1.50E-05|Jy|2009ApJ...698.1682W|typical accuracy|         8 microns   | Broad-band measurement|17 18 44.77 +60 01 15.9 (J2000)| Peak flux|                                        |From reprocessed raw data
24|24 microns (MIPS)   | 1097.299  ||microJy             |1.27E+13|  1.10E-03||Jy|2007ApJ...658..778Y|no uncertainty reported|   23.68   microns   | Broad-band measurement|171844.77 +600115.9 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data; measurementmodified from published value
1|MIPS 24um           | 1.10     |+/-0.33 |milliJy             |1.27E+13|  1.10E-03|+/-0.33E-03 |Jy|1996AJ....111.1431B|uncertainty|1.49       GHz       | Broad-band measurement| | Peak flux|                                        |From new raw data
2|MIPS 70um           | 5.2      |+/-1.7  |milliJy             |4.20E+12|  5.2E-03 |+/-1.7E-03|Jy|2010Natur.464..733S|uncertainty|     71.42 microns   | Broad-band measurement|21 35 11.6 -01 02 52.0 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
25|70 microns (MIPS)   | 5.5       |+/-1.7  | milliJy            |4.20E+12|  5.50E-03|+/-1.70E-03|Jy|2007ApJ...664..713S|estimated error|   71.42   microns   | Broad-band measurement|| Flux in fixed aperture|3 pixel radius aperture                 |From reprocessed raw data
3|MIPS 160um          |          |<30     |milliJy             |1.92E+12|          |30.0E-03|Jy|2009A&A...502..541E|3 sigma|     155.9 microns   | Broad-band measurement| | Flux in fixed aperture|                                        |From reprocessed raw data
4|MAMBO 1200um        | 0.69     |+/-0.54 |milliJy             |2.50E+11|  0.69E-03|+/-0.54E-03|Jy|2004MNRAS.354..779G|uncertainty|      1200 microns   | Broad-band measurement|16 37 06.7 +40 53 15 (J2000)| Flux integrated from map|S/N = 3.81                              |From new raw data
5|VLA 1.4GHz          | 0.34     |+/-0.03 |milliJy             |1.4E9   |  0.34E-3|+/-0.03E-3|Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
28|1.4 GHz (WSRT)      | 0.323     || milliJy            |1.40E+09|  3.23E-04||Jy|2004A&A...424..371M|no uncertainty reported|       1.4 GHz       | Broad-band measurement|17 18 44.781 +60 01 15.14 (J2000)| Flux integrated from map|                                        |From new raw data
29|1.4 GHz (VLA)       | 0.34      ||milliJy             |1.40E+09|  3.40E-04||Jy|2006AJ....131.2859F|no uncertainty reported|     1.4   GHz       | Broad-band measurement|171844.802 +600115.69 (J2000)| Flux integrated from map|                                        |From reprocessed raw data
30|610 MHz (GMRT)      | 0.630     |+/-0.070|milliJy             |6.10E+08|  6.30E-04|+/-7.00E-05|Jy|2007MNRAS.376.1251G|uncertainty|     610   MHz       | Broad-band measurement|17 18 44.83 +60 01 15.8 (J2000)| Flux integrated from map; Pointing corrected|                                        |From new raw data; Corrected for flux in reference beam
