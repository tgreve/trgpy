
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-06-16T05:45:42PDT



Photometric Data for DEEP2 13003805

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|5-10 keV (Chandra)  | 1.59E-15  |+/-0.81E-15|erg/cm^2^/s         |1.81E+18|  8.78E-11|+/-4.48E-11|Jy|2009ApJS..180..102L|1 sigma|      7.50 keV       | Broad-band measurement|214.916980 +52.827245 (J2000)| Modelled datum|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
2|2-10 keV (Chandra)  | 3.89E-15  |+/-0.90E-15|erg/cm^2^/s         |1.45E+18|  2.68E-10|+/-6.21E-11|Jy|2009ApJS..180..102L|1 sigma|      6.00 keV       | Broad-band measurement|214.916980 +52.827245 (J2000)| Modelled datum|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
3|0.5-10 keV (Chandra)| 3.74E-15  |+/-0.62E-15|erg/cm^2^/s         |1.27E+18|  2.94E-10|+/-4.88E-11|Jy|2009ApJS..180..102L|1 sigma|      5.25 keV       | Broad-band measurement|214.916980 +52.827245 (J2000)| Modelled datum|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
4|0.5-2 keV (Chandra) | 0.70E-15  |+/-0.18E-15|erg/cm^2^/s         |3.02E+17|  2.32E-10|+/-5.96E-11|Jy|2009ApJS..180..102L|1 sigma|      1.25 keV       | Broad-band measurement|214.916980 +52.827245 (J2000)| Modelled datum|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
5|CO(3-2) (PdBI)      ||<0.15      |Jy km/s             |3.46E+11|  1.16E+06|7.76E+04|Jy-Hz|2010Natur.463..781T|3 sigma|   345.998 GHz       | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|                                        |From new raw data
