
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-07-08T03:43:25PDT



Photometric Data for SDSS J123646.20+621142.4

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|U_300 (WFPC-2)      | 23.21     ||mag                 |1.02E+15|  5.36E-07||Jy|1996AJ....112.1335W|no uncertainty reported|2942       A         | Broad-band measurement|123646.20 +621141.2 (J2000)| Flux integrated from map|                                        |From new raw data; derived from a flux in a different bandand a color
2|U_300_ (HST)        | 1610.00   |+/-32.31|nJy                 |1.02E+15|  1.61E-06|+/-3.23E-08|Jy|1999ApJ...513...34F|1 sigma|2942       A         | Broad-band measurement|| Flux in fixed aperture|                                        |From reprocessed raw data
3|U (KPNO) AB         | 23.2      || mag                |8.22E+14|  1.91E-06||Jy|2004AJ....127.3137C|no uncertainty reported| 3647.65   A         | Broad-band measurement|189.192429 +62.19511 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
4|B F435W (HST/ACS) AB      | 22.802    ||mag                 |6.98E+14|  2.75E-06||Jy|2007ApJ...660...81M|no uncertainty reported|    4297   A         | Broad-band measurement|12 36 46.189 +62 11 41.97 (J2000)| Flux integrated from map|                                        |From reprocessed raw data; Corrected for contaminatingsources
5|B (Subaru) AB       | 23.14     ||mag                 |6.77E+14|  2.01E-06||Jy|2006ApJ...653.1027W|no uncertainty reported| 4427.60   A         | Broad-band measurement|189.192454 62.194992 (J2000)| Flux in fixed aperture|3" diameter aperture                    |Averaged from previously published data
6|B (Subaru) AB       | 23.2      || mag                |6.77E+14|  1.91E-06||Jy|2004AJ....127.3137C|no uncertainty reported| 4427.60   A         | Broad-band measurement|189.192429 +62.19511 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
7|B_450 (WFPC-2)      | 22.71     ||mag                 |6.63E+14|  3.59E-06||Jy|1996AJ....112.1335W|no uncertainty reported|4519       A         | Broad-band measurement|123646.20 +621141.2 (J2000)| Flux integrated from map|                                        |From new raw data; derived from a flux in a different bandand a color
8|B_450_ (HST)        | 2679.00   |+/-15.73|nJy                 |6.63E+14|  2.68E-06|+/-1.57E-08|Jy|1999ApJ...513...34F|1 sigma|4519       A         | Broad-band measurement|| Flux in fixed aperture|                                        |From reprocessed raw data
9|V (Subaru) AB       | 22.8      || mag                |5.48E+14|  2.75E-06||Jy|2004AJ....127.3137C|no uncertainty reported| 5471.22   A         | Broad-band measurement|189.192429 +62.19511 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
10|V (HST/ACS) AB      | 22.169    ||mag                 |5.08E+14|  4.93E-06||Jy|2007ApJ...660...81M|no uncertainty reported|    5907   A         | Broad-band measurement|12 36 46.189 +62 11 41.97 (J2000)| Flux integrated from map|                                        |From reprocessed raw data; Corrected for contaminatingsources
11|V_606_ (HST)        | 4358.00   |+/-11.40|nJy                 |5.05E+14|  4.36E-06|+/-1.14E-08|Jy|1999ApJ...513...34F|1 sigma|5934       A         | Broad-band measurement|| Flux in fixed aperture|                                        |From reprocessed raw data
12|V_606 (WFPC-2)      | 22.18     ||mag                 |5.05E+14|  4.57E-06||Jy|1996AJ....112.1335W|no uncertainty reported|5934       A         | Broad-band measurement|123646.20 +621141.2 (J2000)| Flux integrated from map|                                        |From new raw data
13|R (Keck II) AB      | 22.25     || mag                |4.62E+14|  4.57E-06||Jy|2004AJ....127.3121W|no uncertainty reported|   648.7   A         | Broad-band measurement|12 36 46.189 +62 11 41.97 (J2000)| Total flux|                                        |From new raw data
14|R (Subaru) AB       | 22.30     ||mag                 |4.59E+14|  4.37E-06||Jy|2006ApJ...653.1027W|no uncertainty reported| 6534.16   A         | Broad-band measurement|189.192454 62.194992 (J2000)| Flux in fixed aperture|3" diameter aperture                    |Averaged from previously published data
15|R (Subaru) AB       | 22.3      || mag                |4.59E+14|  4.37E-06||Jy|2004AJ....127.3137C|no uncertainty reported| 6534.16   A         | Broad-band measurement|189.192429 +62.19511 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
16|i F775W (HST/ACS) AB      | 21.400    ||mag                 |3.86E+14|  1.00E-05||Jy|2007ApJ...660...81M|no uncertainty reported|    7764   A         | Broad-band measurement|12 36 46.189 +62 11 41.97 (J2000)| Flux integrated from map|                                        |From reprocessed raw data; Corrected for contaminatingsources
17|I_814 (WFPC-2)      | 21.23     ||mag                 |3.78E+14|  8.02E-06||Jy|1996AJ....112.1335W|no uncertainty reported|7924       A         | Broad-band measurement|123646.20 +621141.2 (J2000)| Flux integrated from map|                                        |From new raw data; derived from a flux in a different bandand a color
18|I_814_ (HST)        | 10710.00  |+/-20.51|nJy                 |3.78E+14|  1.07E-05|+/-2.05E-08|Jy|1999ApJ...513...34F|1 sigma|7924       A         | Broad-band measurement|| Flux in fixed aperture|                                        |From reprocessed raw data
19|AB(814) Best        | 21.26     ||mag                 |3.78E+14|  1.14E-05||Jy|1999ApJ...513...34F|no uncertainty reported| 7924      A         | Broad-band measurement|123646.166 +621142.09 (     )| Flux in fixed aperture|                                        |From reprocessed raw data; Corrected for contaminatingsources
20|I (Subaru) AB       | 21.6      || mag                |3.76E+14|  8.32E-06||Jy|2004AJ....127.3137C|no uncertainty reported| 7975.89   A         | Broad-band measurement|189.192429 +62.19511 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
21|I (Subaru) AB       | 21.59     ||mag                 |3.76E+14|  8.40E-06||Jy|2006ApJ...653.1027W|no uncertainty reported| 7975.89   A         | Broad-band measurement|189.192454 62.194992 (J2000)| Flux in fixed aperture|3" diameter aperture                    |Averaged from previously published data
22|F814W (HST) AB      | 21.30     ||mag                 |3.60E+14|  1.10E-05||Jy|2004AJ....127..131S|no uncertainty reported|    8333   A         | Broad-band measurement|12 36 46.18 +62 11 42.1 (J2000)| Flux in fixed aperture|                                        |From new raw data; derived from a flux in a different bandand a color
23|z' (Subaru) AB      | 21.2      || mag                |3.31E+14|  1.20E-05||Jy|2004AJ....127.3137C|no uncertainty reported| 9069.21   A         | Broad-band measurement|189.192429 +62.19511 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
24|z F850LP (HST/ACS) AB      | 20.776    ||mag                 |3.17E+14|  1.78E-05||Jy|2007ApJ...660...81M|no uncertainty reported|    9445   A         | Broad-band measurement|12 36 46.189 +62 11 41.97 (J2000)| Flux integrated from map|                                        |From reprocessed raw data; Corrected for contaminatingsources
25|J (KPNO)            | 33010.    |+/-497. |nJy                 |2.38E+14|  3.30E-05|+/-4.97E-07|Jy|1999ApJ...513...34F|1 sigma|1.26       microns   | Broad-band measurement|| Flux in fixed aperture|                                        |From reprocessed raw data
26|H (KPNO)            | 43280.    |+/-883. |nJy                 |1.87E+14|  4.33E-05|+/-8.83E-07|Jy|1999ApJ...513...34F|1 sigma|1.60       microns   | Broad-band measurement|| Flux in fixed aperture|                                        |From reprocessed raw data
27|F160W (HST) AB      | 19.88     ||mag                 |1.86E+14|  4.06E-05||Jy|2004AJ....127..131S|no uncertainty reported|   1.608   microns   | Broad-band measurement|12 36 46.18 +62 11 42.1 (J2000)| Total flux|                                        |From new raw data
28|HK' (UH) AB         | 19.9      || mag                |1.58E+14|  3.98E-05||Jy|2004AJ....127.3137C|no uncertainty reported|18947.38   A         | Broad-band measurement|189.192429 +62.19511 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
29|HK' (QUIRC) AB      | 19.88     |+/-0.03 |mag                 |1.58E+14|  4.06E-05|+/-1.12E-06|Jy|2006ApJ...653.1027W|uncertainty|18947.38   A         | Broad-band measurement|189.192454 62.194992 (J2000)| Flux in fixed aperture|3" diameter aperture                    |Averaged from previously published data
30|K (KPNO)            | 66470.    |+/-786. |nJy                 |1.35E+14|  6.65E-05|+/-7.86E-07|Jy|1999ApJ...513...34F|1 sigma|2.22       microns   | Broad-band measurement|| Flux in fixed aperture|                                        |From reprocessed raw data
31|3.6 microns (IRAC)  | 97.70     |+/-4.89 |microJy             |8.44E+13|  9.77E-05|+/-4.89E-06|Jy|2011AJ....141....1T|rms uncertainty|     3.550 microns   | Broad-band measurement|189.192490 62.195011 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
32|4.5 microns (IRAC)  | 72.60     |+/-3.63 |microJy             |6.67E+13|  7.26E-05|+/-3.63E-06|Jy|2011AJ....141....1T|rms uncertainty|     4.493 microns   | Broad-band measurement|189.192490 62.195011 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
33|5.8 microns (IRAC)  | 52.20     |+/-2.64 |microJy             |5.23E+13|  5.22E-05|+/-2.64E-06|Jy|2011AJ....141....1T|rms uncertainty|     5.731 microns   | Broad-band measurement|189.192490 62.195011 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
34|8.0 microns (IRAC)  | 44.60     |+/-2.28 |microJy             |3.81E+13|  4.46E-05|+/-2.28E-06|Jy|2011AJ....141....1T|rms uncertainty|     7.872 microns   | Broad-band measurement|189.192490 62.195011 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
35|11 microns (AKARI)  | 61.0      |+/-15   | microJy            |2.73E+13|  6.10E-05|+/-1.50E-05|Jy|2009MNRAS.394..375N|uncertainty|        11 microns   | Broad-band measurement|12 36 46.18 +62 11 42.41 (J2000)| Flux integrated from map|                                        |From new raw data
36|15 microns (ISOCAM) | 125       |+/-41   |microJy             |2.00E+13|  1.25E-04|+/-4.10E-05|Jy|2006A&A...451...57M|68% confidence|    15.0   microns   | Broad-band measurement|189.1924133 62.1951141 (J2000)| Flux integrated from map|                                        |Averaged from previously published data
37|16 microns (IRS)    | 245.7     |+/-11.7 |microJy             |1.90E+13|  2.46E-04|+/-1.17E-05|Jy|2011AJ....141....1T|rms uncertainty|      15.8 microns   | Broad-band measurement|189.192490 62.195011 (J2000)| From fitting to map|                                        |From new raw data
38|16 microns (IRS)    | 275       |+/-18   | microJy            |1.87E+13|  2.75E-04|+/-1.80E-05|Jy|2009MNRAS.394..375N|uncertainty|        16 microns   | Broad-band measurement|12 36 46.18 +62 11 42.41 (J2000)| Flux integrated from map|                                        |Averaged from previously published data
39|18 microns (AKARI)  | 212       |+/-37   | microJy            |1.67E+13|  2.12E-04|+/-3.70E-05|Jy|2009MNRAS.394..375N|uncertainty|        18 microns   | Broad-band measurement|12 36 46.18 +62 11 42.41 (J2000)| Flux integrated from map|                                        |From new raw data
40|24 microns (MIPS)   | 290       |+/-5    |microJy             |1.27E+13|  2.90E-04|+/-5.00E-06|Jy|2006A&A...451...57M|68% confidence|   23.68   microns   | Broad-band measurement|189.1924133 62.1951141 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
41|24 microns (MIPS)   | 293.0     |+/-5.5  |microJy             |1.27E+13|  2.93E-04|+/-5.50E-06|Jy|2011AJ....141....1T|rms uncertainty|     23.68 microns   | Broad-band measurement|189.192490 62.195011 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
42|24 microns (MIPS)   | 299.1     |+/-2.5  |microJy             |1.27E+13|  2.99E-04|+/-2.50E-06|Jy|2011A&A...528A..35M|uncertainty|     23.68 microns   | Broad-band measurement|12 36 46.20 +62 11 41.97 (J2000)| Flux integrated from map|                                        |From new raw data
1|MIPS 24 microns      | 300.      |+/-6.0  |microJy         |1.25E+13 |  300.E-06|+/-6.0E-06  |Jy |1990IRASF.C...0000M|3sigma uncertainty| 25        microns   | Broad-band measurement|115813.1 +302058 (B1950)| Flux in fixed aperture|                                        |From new raw data
43|70 microns (MIPS)   ||<3.1       |milliJy             |4.20E+12||3.10E-03|Jy|2011A&A...528A..35M|no uncertainty reported|     71.42 microns   | Broad-band measurement|12 36 46.20 +62 11 41.97 (J2000)| Flux integrated from map|                                        |From new raw data
2|70 microns (PACS)    |           |<2.0    |mJy             |4.283e+12|          |2.0E-03     |Jy |2.40e+01           |3sigma |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
3|100 microns (PACS)   | 2.9       |+/-0.3  |mJy             |2.998e+12|  2.9E-03 |+/-0.3E-03  |Jy |2.40e+01           |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
4|160 microns (PACS)   | 5.8       |+/-0.7  |mJy             |1.874e+12|  5.8E-03 |+/-0.7E-03  |Jy |2.40e+01           |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
5|250 microns (SPIRE)  | 12.7      |+/-2.5  |mJy             |1.199e+12|  12.7E-03|+/-2.5e-03  |Jy |2.40e+01           |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
6|350 microns (SPIRE)  | 10.7      |+/-3.0  |mJy             |8.565e+11|  10.7E-03|+/-3.0e-03  |Jy |2.40e+01           |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
7|500 microns (SPIRE)  |           |<12.0   |mJy             |5.996e+11|          |12.0e-03    |Jy |2.40e+01           |3sigma |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
8|1160 microns (Penner)|           |<1.7    |mJy             |2.58442E+11|        |1.7E-03     |Jy |2004MNRAS.354..779G|3sigma uncertainty|      1200 microns   | Broad-band measurement|16 36 55.9 +40 59 12 (J2000)| Flux integrated from map|S/N = 3.66                              |From new raw data
44|1.4 GHz (VLA)       | 21.04     ||microJy             |1.40E+09|  2.10E-05||Jy|2006A&A...451...57M|no uncertainty reported|     1.4   GHz       | Broad-band measurement|189.1924133 62.1951141 (J2000)| Flux integrated from map|                                        |From new raw data
