
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-07-08T05:21:33PDT



Photometric Data for GOODS J123750.89+621601.1

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|4.0-8 keV (Chandra) ||<0.85E-15  |ergs cm^-2^ s^-1^   |1.45E+18||5.86E-11|Jy|2003AJ....126..539A|3 sigma|       6   keV       | Broad-band measurement|12 37 50.88 +62 16 01.0 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
2|2.0-8 keV (Chandra) ||<0.63E-15  |ergs cm^-2^ s^-1^   |1.21E+18||5.21E-11|Jy|2003AJ....126..539A|3 sigma|       5   keV       | Broad-band measurement|12 37 50.88 +62 16 01.0 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
3|0.5-8 keV (Chandra) | 0.69E-15  ||ergs cm^-2^ s^-1^   |1.03E+18|  6.71E-11||Jy|2003AJ....126..539A|no uncertainty reported|    4.25   keV       | Broad-band measurement|12 37 50.88 +62 16 01.0 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
4|2.0-4 keV (Chandra) ||<0.21E-15  |ergs cm^-2^ s^-1^   |7.25E+17||2.89E-11|Jy|2003AJ....126..539A|3 sigma|       3   keV       | Broad-band measurement|12 37 50.88 +62 16 01.0 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
5|1.0-2 keV (Chandra) | 0.07E-15  ||ergs cm^-2^ s^-1^   |3.63E+17|  1.93E-11||Jy|2003AJ....126..539A|no uncertainty reported|     1.5   keV       | Broad-band measurement|12 37 50.88 +62 16 01.0 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
6|0.5-2 keV (Chandra) | 0.10E-15  ||ergs cm^-2^ s^-1^   |3.02E+17|  3.31E-11||Jy|2003AJ....126..539A|no uncertainty reported|    1.25   keV       | Broad-band measurement|12 37 50.88 +62 16 01.0 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
7|0.5-1 keV (Chandra) ||<0.07E-15  |ergs cm^-2^ s^-1^   |1.81E+17||3.86E-11|Jy|2003AJ....126..539A|3 sigma|    0.75   keV       | Broad-band measurement|12 37 50.88 +62 16 01.0 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
8|U (KPNO) AB         | 24.7      || mag                |8.22E+14|  4.79E-07||Jy|2004AJ....127.3137C|no uncertainty reported| 3647.65   A         | Broad-band measurement|189.462051 +62.26698 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
9|F435W (HST) AB      | 21.007    |+/-0.006|mag                 |6.92E+14|  1.44E-05|+/-7.94E-08|Jy|2011ApJ...734..121S|uncertainty|      4333 A         | Broad-band measurement|189.462021 62.266979 (J2000)| Total flux|                                        |From reprocessed raw data
10|F435W (HST) AB      | 21.07     |+/-0.21 |mag                 |6.92E+14|  1.36E-05|+/-2.62E-06|Jy|2011ApJ...734..121S|uncertainty|      4333 A         | Broad-band measurement|189.462021 62.266979 (J2000)| Modelled datum|Host galaxy mag                         |From reprocessed raw data
11|F435W (HST) AB      | 24.12     |+/-0.14 |mag                 |6.92E+14|  8.17E-07|+/-1.05E-07|Jy|2011ApJ...734..121S|uncertainty|      4333 A         | Broad-band measurement|189.462021 62.266979 (J2000)| Modelled datum|Central point source mag                |From reprocessed raw data
12|B (Subaru) AB       | 24.4      || mag                |6.77E+14|  6.31E-07||Jy|2004AJ....127.3137C|no uncertainty reported| 4427.60   A         | Broad-band measurement|189.462051 +62.26698 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
13|V (Subaru) AB       | 23.9      || mag                |5.48E+14|  1.00E-06||Jy|2004AJ....127.3137C|no uncertainty reported| 5471.22   A         | Broad-band measurement|189.462051 +62.26698 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
14|R (Keck II) AB      | 22.99     || mag                |4.62E+14|  2.31E-06||Jy|2004AJ....127.3121W|no uncertainty reported|   648.7   A         | Broad-band measurement|12 37 50.887 +62 16 00.69 (J2000)| Total flux|                                        |From new raw data
15|R (Subaru) AB       | 23.0      || mag                |4.59E+14|  2.29E-06||Jy|2004AJ....127.3137C|no uncertainty reported| 6534.16   A         | Broad-band measurement|189.462051 +62.26698 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
16|I (Subaru) AB       | 22.1      || mag                |3.76E+14|  5.25E-06||Jy|2004AJ....127.3137C|no uncertainty reported| 7975.89   A         | Broad-band measurement|189.462051 +62.26698 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
17|z' (Subaru) AB      | 21.3      || mag                |3.31E+14|  1.10E-05||Jy|2004AJ....127.3137C|no uncertainty reported| 9069.21   A         | Broad-band measurement|189.462051 +62.26698 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
18|HK' (UH) AB         | 19.6      || mag                |1.58E+14|  5.25E-05||Jy|2004AJ....127.3137C|no uncertainty reported|18947.38   A         | Broad-band measurement|189.462051 +62.26698 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
19|3.6 microns (IRAC)  | 119.00    |+/-5.95 |microJy             |8.44E+13|  1.19E-04|+/-5.95E-06|Jy|2011AJ....141....1T|rms uncertainty|     3.550 microns   | Broad-band measurement|189.462051 62.266884 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
20|4.5 microns (IRAC)  | 98.60     |+/-4.93 |microJy             |6.67E+13|  9.86E-05|+/-4.93E-06|Jy|2011AJ....141....1T|rms uncertainty|     4.493 microns   | Broad-band measurement|189.462051 62.266884 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
21|5.8 microns (IRAC)  | 65.40     |+/-3.30 |microJy             |5.23E+13|  6.54E-05|+/-3.30E-06|Jy|2011AJ....141....1T|rms uncertainty|     5.731 microns   | Broad-band measurement|189.462051 62.266884 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
22|8.0 microns (IRAC)  | 53.50     |+/-2.72 |microJy             |3.81E+13|  5.35E-05|+/-2.72E-06|Jy|2011AJ....141....1T|rms uncertainty|     7.872 microns   | Broad-band measurement|189.462051 62.266884 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
23|16 microns (IRS)    | 164.5     |+/-11.8 |microJy             |1.90E+13|  1.65E-04|+/-1.18E-05|Jy|2011AJ....141....1T|rms uncertainty|      15.8 microns   | Broad-band measurement|189.462051 62.266884 (J2000)| From fitting to map|                                        |From new raw data
24|24 microns (MIPS)   | 186.0     |+/-5.4  |microJy             |1.27E+13|  1.86E-04|+/-5.40E-06|Jy|2011AJ....141....1T|rms uncertainty|     23.68 microns   | Broad-band measurement|189.462051 62.266884 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
25|24 microns (MIPS)   | 191.4     |+/-2.6  |microJy             |1.27E+13|  1.91E-04|+/-2.60E-06|Jy|2011A&A...528A..35M|uncertainty|     23.68 microns   | Broad-band measurement|12 37 50.89 +62 16 00.71 (J2000)| Flux integrated from map|                                        |From new raw data
1|MIPS 24 microns      | 188.    |+/-6.0 |microJy         |1.25E+13 |  188.E-06|+/-6.0E-06 |Jy|1990IRASF.C...0000M|3sigma uncertainty| 25        microns   | Broad-band measurement|115813.1 +302058 (B1950)| Flux in fixed aperture|                                        |From new raw data
2|70 microns (PACS)    |         |<2.0   |mJy             |4.283e+12|          |2.0E-03 |Jy |2.40e+01 |3sigma |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
26|70 microns (MIPS)   ||<2.4       |milliJy             |4.20E+12||2.40E-03|Jy|2011A&A...528A..35M|no uncertainty reported|     71.42 microns   | Broad-band measurement|12 37 50.89 +62 16 00.71 (J2000)| Flux integrated from map|                                        |From new raw data
3|100 microns (PACS)   | 1.7     |+/-0.3 |mJy             |2.998e+12|  1.7E-03 |+/-0.3E-03 |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
4|160 microns (PACS)   | 4.8     |+/-1.1 |mJy             |1.874e+12|  4.8E-03 |+/-1.1E-03 |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
5|250 microns (SPIRE)  | 8.6     |+/-2.5 |mJy             |1.199e+12|  8.6E-03 |+/-2.5e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
6|350 microns (SPIRE)  | 8.8     |+/-3.0 |mJy             |8.565e+11|  8.8E-03 |+/-3.0e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
7|500 microns (SPIRE)  |         |<12.0  |mJy             |5.996e+11|          |12.0e-03  |Jy |2.40e+01 |3sigma |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
8|1160 microns (Penner)|         |<1.8   |mJy             |2.58442E+11|        |1.8E-03|Jy|2004MNRAS.354..779G|3sigma uncertainty|      1200 microns   | Broad-band measurement|16 36 55.9 +40 59 12 (J2000)| Flux integrated from map|S/N = 3.66                              |From new raw data
27|1.4 GHz (VLA)       | 27.7      |+/-5.7  |microJy             |1.40E+09|  2.77E-05|+/-5.70E-06|Jy|2010ApJS..188..178M|uncertainty|       1.4 GHz       | Broad-band measurement|12 37 50.84 +62 16 00.7 (J2000)| Total flux; Beam filling or dilution corrected|Major=1.4"; Minor=0.0"; PA=114 deg      |From new raw data
