
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-07-08T05:55:10PDT



Photometric Data for GNS 0856

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|U (KPNO) AB         | 28.94     ||mag                 |8.44E+14|  9.64E-09||Jy|2006ApJ...653.1004R|no uncertainty reported|    3550   A         | Broad-band measurement|123642.96 +620958.1 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data; derived from aflux in a different band and a color
2|G (KECK) AB         | 26.48     ||mag                 |6.27E+14|  9.29E-08||Jy|2006ApJ...653.1004R|no uncertainty reported|    4780   A         | Broad-band measurement|123642.96 +620958.1 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data; derived from aflux in a different band and a color
3|R (KECK) AB         | 25.48     ||mag                 |4.39E+14|  2.33E-07||Jy|2006ApJ...653.1004R|no uncertainty reported|    6830   A         | Broad-band measurement|123642.96 +620958.1 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data
8|I (Cousins)         | 25.9     |+/-0.1 |mag           |3.79E+14|  999.E-01|+/-99.E-03|Jy|Add flux in Jy|1 sigma|    7900   A         | Broad-band measurement| | Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
4|J (WIRC) AB         | 22.86     ||mag                 |2.40E+14|  2.61E-06||Jy|2006ApJ...653.1004R|no uncertainty reported|   1.250   microns   | Broad-band measurement|123642.96 +620958.1 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data
5|F160W (HST) AB      | 21.77     |+/-0.05 |mag                 |1.87E+14|  7.11E-06|+/-3.27E-07|Jy|2011MNRAS.413...80C|uncertainty|      1.60 microns   | Broad-band measurement|189.178649 62.166355 (J2000)| Total flux|                                        |From new raw data
6|K_s (WIRC) AB       | 21.04     ||mag                 |1.39E+14|  1.39E-05||Jy|2006ApJ...653.1004R|no uncertainty reported|   2.150   microns   | Broad-band measurement|123642.96 +620958.1 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data
7|3.6 microns IRAC AB | 20.59     |+/-0.07 |mag                 |8.44E+13|  2.11E-05|+/-1.36E-06|Jy|2006ApJ...653.1004R|uncertainty|   3.550   microns   | Broad-band measurement|123642.96 +620958.1 (J2000)| Flux integrated from map|                                        |From new raw data
8|4.5 microns IRAC AB | 20.50     |+/-0.07 |mag                 |6.67E+13|  2.29E-05|+/-1.48E-06|Jy|2006ApJ...653.1004R|uncertainty|   4.493   microns   | Broad-band measurement|123642.96 +620958.1 (J2000)| Flux integrated from map|                                        |From new raw data
9|5.8 microns IRAC AB | 20.33     |+/-0.07 |mag                 |5.23E+13|  2.68E-05|+/-1.73E-06|Jy|2006ApJ...653.1004R|uncertainty|   5.731   microns   | Broad-band measurement|123642.96 +620958.1 (J2000)| Flux integrated from map|                                        |From new raw data
10|8.0 microns IRAC AB | 20.76     |+/-0.08 |mag                 |3.81E+13|  1.80E-05|+/-1.33E-06|Jy|2006ApJ...653.1004R|uncertainty|   7.872   microns   | Broad-band measurement|123642.96 +620958.1 (J2000)| Flux integrated from map|                                        |From new raw data
11|24 microns (MIPS)   | 21.0      |+/-4.8  |microJy             |1.27E+13|  2.10E-05|+/-4.80E-06|Jy|2006ApJ...653.1004R|uncertainty|   23.68   microns   | Broad-band measurement|123642.96 +620958.1 (J2000)| Flux integrated from map|                                        |From new raw data
34|24 microns (MIPS)   |      |<15  |microJy             |1.27E+13|  |15.0E-06|Jy|2011AJ....141....1T|3sigma uncertainty|     23.68 microns   | Broad-band measurement|189.300690 62.298355 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
36|70 microns (MIPS)   ||<1.9       |milliJy             |4.20E+12||1.9E-03|Jy|2011A&A...528A..35M|3sigma uncertainty reported|     71.42 microns   | Broad-band measurement|12 37 12.17 +62 17 54.01 (J2000)| Flux integrated from map|                                        |From new raw data
29|850 microns (SCUBA) |        |<3.4  |milliJy             |3.53E+11|  |3.40E-03|Jy|2005ApJ...622..772C|3sigma uncertainty|     850   microns   | Broad-band measurement|123600.15 +621047.2 (J2000)| Flux integrated from map|                                        |From new raw data
7|1200 microns (MAMBO)|           |<0.9    |mJy                 |2.50E+11|          |0.9E-03|Jy|2004MNRAS.354..779G|3sigma uncertainty|      1200 microns   | Broad-band measurement|16 36 55.9 +40 59 12 (J2000)| Flux integrated from map|S/N = 3.66                              |From new raw data
12|1.4 GHz (VLA)       | 24.0      |+/-4.3  |microJy             |1.40E+09|  2.40E-05|+/-4.30E-06|Jy|2010ApJS..188..178M|uncertainty|       1.4 GHz       | Broad-band measurement|12 36 42.86 +62 09 58.5 (J2000)| Total flux; Beam filling or dilution corrected|Major=0.0"; Minor=0.0"; PA=0 deg        |From new raw data
