
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-02-19T12:06:08PST


z=2.4494
Photometric Data for SMM J163658.19+410523.8

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
6|I (Cousins)         | 24.48     |+/-0.20 |mag                 |3.79E+14|  4.12E-07|+/-8.33E-08|Jy|2004ApJ...616...71S|1 sigma|    7900   A         | Broad-band measurement| | Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
6|F160W (HST/NICMOS)  | 24.41    |+/-0.08| mag                |1.87E+14|  6.25173e-07|+/-4.6064425e-08|Jy|2007A&A...470..467C|internal error|       1.6 microns   | Broad-band measurement| | From fitting to map|                                        |From new raw data
11|K_s_ (2MASS)        | 19.77     |+/-0.06 |mag                 |1.38E+14|  8.24E-06|+/-4.68E-07|Jy|2004ApJ...616...71S|1 sigma|    2.17   microns   | Broad-band measurement| | Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
12|K (GeminiN)         | 20.77     |+/-0.27 |mag                 |1.36E+14|  3.15E-06|+/-7.83E-07|Jy|2011MNRAS.412..295T|uncertainty|      2.21 microns   | Broad-band measurement|| Flux in fixed aperture|6" diameter aperture                    |From new raw data
13|3.6 microns (IRAC)  | 1.9588E+01|+/-2.2813E-01|microJy             |8.44E+13|  1.96E-05|+/-2.28E-07|Jy|2013SSTSLC4.2....0C|uncertainty|3.55       microns   | Broad-band measurement|| Flux in fixed aperture|5.8" aperture                           |From new raw data
14|3.6 microns (IRAC)  | 1.5518E+01|+/-1.7771E-01|microJy             |8.44E+13|  1.55E-05|+/-1.78E-07|Jy|2013SSTSLC4.2....0C|uncertainty|3.55       microns   | Broad-band measurement|| Flux in fixed aperture|3.8" aperture                           |From new raw data
12|3.6 microns (IRAC)  | 15.3      |+/-1.6  |microJy             |8.44E+13|  1.53E-05|+/-1.60E-06|Jy|2009ApJ...699.1610H|uncertainty|     3.550 microns   | Broad-band measurement|16 36 58.13 +41 05 23.1 (J2000)| Flux in fixed aperture|                                        |From new raw data
16|4.5 microns (IRAC)  | 2.1366E+01|+/-2.7777E-01|microJy             |6.67E+13|  2.14E-05|+/-2.78E-07|Jy|2013SSTSLC4.2....0C|uncertainty|4.493      microns   | Broad-band measurement|| Flux in fixed aperture|3.8" aperture                           |From new raw data
17|4.5 microns (IRAC)  | 2.5335E+01|+/-3.8407E-01|microJy             |6.67E+13|  2.53E-05|+/-3.84E-07|Jy|2013SSTSLC4.2....0C|uncertainty|4.493      microns   | Broad-band measurement|| Flux in fixed aperture|5.8" aperture                           |From new raw data
13|4.5 microns (IRAC)  | 21.8      |+/-2.4  |microJy             |6.67E+13|  2.18E-05|+/-2.40E-06|Jy|2009ApJ...699.1610H|uncertainty|     4.493 microns   | Broad-band measurement|16 36 58.13 +41 05 23.1 (J2000)| Flux in fixed aperture|                                        |From new raw data
19|5.8 microns (IRAC)  | 2.8592E+01|+/-1.3293E+00|microJy             |5.23E+13|  2.86E-05|+/-1.33E-06|Jy|2013SSTSLC4.2....0C|uncertainty|5.731      microns   | Broad-band measurement|| Flux in fixed aperture|3.8" aperture                           |From new raw data
20|5.8 microns (IRAC)  | 3.6898E+01|+/-1.8417E+00|microJy             |5.23E+13|  3.69E-05|+/-1.84E-06|Jy|2013SSTSLC4.2....0C|uncertainty|5.731      microns   | Broad-band measurement|| Flux in fixed aperture|5.8" aperture                           |From new raw data
14|5.8 microns (IRAC)  | 28.9      |+/-3.2  |microJy             |5.23E+13|  2.89E-05|+/-3.20E-06|Jy|2009ApJ...699.1610H|uncertainty|     5.731 microns   | Broad-band measurement|16 36 58.13 +41 05 23.1 (J2000)| Flux in fixed aperture|                                        |From new raw data
23|8.0 microns (IRAC)  | 3.4146E+01|+/-2.4287E+00|microJy             |3.81E+13|  3.41E-05|+/-2.43E-06|Jy|2013SSTSLC4.2....0C|uncertainty|7.872      microns   | Broad-band measurement|| Flux in fixed aperture|5.8" aperture                           |From new raw data
24|8.0 microns (IRAC)  | 3.3253E+01|+/-1.8145E+00|microJy             |3.81E+13|  3.33E-05|+/-1.81E-06|Jy|2013SSTSLC4.2....0C|uncertainty|7.872      microns   | Broad-band measurement|| Flux in fixed aperture|3.8" aperture                           |From new raw data
15|8.0 microns (IRAC)  | 29.9      |+/-3.5  |microJy             |3.85E+13|  2.99E-05|+/-3.50E-06|Jy|2009ApJ...699.1610H|uncertainty|     7.782 microns   | Broad-band measurement|16 36 58.13 +41 05 23.1 (J2000)| Flux in fixed aperture|                                        |From new raw data
16|24 microns (MIPS)   | 330.0     |+/-55.0 |microJy             |1.27E+13|  3.30E-04|+/-5.50E-05|Jy|2009ApJ...699.1610H|uncertainty|     23.68 microns   | Broad-band measurement|163658.19 +410523.8 (J2000)| Flux in fixed aperture|                                        |From new raw data
17|24 microns (Spitzer)| 330       |+/-55   |microJy             |1.27E+13|  3.30E-04|+/-5.50E-05|Jy|2011ApJ...726...93R|uncertainty|     23.68 microns   | Broad-band measurement|16 36 58.19 +41 05 23.8 (J2000)| Not reported in paper|                                        |Averaged from previously published data
27|24 microns (MIPS)   | 3.9549E+02|+/-3.8397E+01|microJy             |1.27E+13|  3.95E-04|+/-3.84E-05|Jy|2013SSTSLC4.2....0C|uncertainty|23.68      microns   | Broad-band measurement|| Modelled datum|PSF fit                                 |From new raw data
28|24 microns (MIPS)   | 5.4406E+02|+/-3.5605E+01|microJy             |1.27E+13|  5.44E-04|+/-3.56E-05|Jy|2013SSTSLC4.2....0C|uncertainty|23.68      microns   | Broad-band measurement|| Flux in fixed aperture|14.7" aperture                          |From new raw data
18|70 microns (MIPS)   | |<7.9       |milliJy             |4.20E+12| |7.90E-03|Jy|2009ApJ...699.1610H|3 sigma|     71.42 microns   | Broad-band measurement|163658.19 +410523.8 (J2000)| Flux in fixed aperture|                                        |From new raw data
19|350 microns (SHARC2)| 45.2      |+/-5.3  |milliJy             |8.57E+11|  4.52E-02|+/-5.30E-03|Jy|2006ApJ...650..592K|uncertainty|     350   microns   | Broad-band measurement| | Total flux|                                        |From new raw data
21|850 microns (SCUBA) | 10.7      |+/-2.0  |milliJy             |3.53E+11|  1.07E-02|+/-2.00E-03|Jy|2005ApJ...622..772C|uncertainty|     850   microns   | Broad-band measurement|163658.19 +410523.8 (J2000)| Flux integrated from map|                                        |From new raw data
22|850 microns (SCUBA) | 11.0      |+/-1.9  |mag                 |3.53E+11|  1.10E-02|+/-1.90E-03|Jy|2006MNRAS.370.1057S|uncertainty|     850   microns   | Broad-band measurement|16 36 58.62 +41 05 24.9 (J2000)| From fitting to map|S/N = 6.92                              |From reprocessed raw data
28|234.456 GHz (PdBI)  | 2.0       |+/-0.2  |milliJy             |2.34E+11|  2.00E-03|+/-2.00E-04|Jy|2011ApJ...730...18W|uncertainty|   234.456 GHz       | Broad-band measurement|16 36 58.17 +41 05 23.3 (J2000)| Flux integrated from map|                                        |From new raw data
25|1.3 mm (PdBI)       | 1.5       |+/-0.5  |milliJy             |2.31E+11|  1.50E-03|+/-5.00E-04|Jy|2006ApJ...640..228T|uncertainty|     1.3   mm        | Broad-band measurement| | Flux integrated from map|                                        |From new raw data
30|142.573 GHz (PdBI)  | 0.6       ||milliJy             |1.43E+11|  6.00E-04||Jy|2011ApJ...730...18W|no uncertainty reported|   142.573 GHz       | Broad-band measurement|16 36 58.17 +41 05 23.3 (J2000)| Flux integrated from map|                                        |From new raw data
26|1.4 GHz (VLA)       | 97        |+/-11   | microJy            |1.40E+09|  9.70E-05|+/-1.10E-05|Jy|2006MNRAS.371..963B|1 sigma|       1.4 GHz       | Broad-band measurement|16 36 58.179 +41 05 23.78 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
27|1.4 GHz (VLA)       | 115        |+/-11   | microJy            |1.40E+09|  11.5E-05|+/-1.10E-05|Jy|2006MNRAS.371..963B|1 sigma|       1.4 GHz       | Broad-band measurement|16 36 58.179 +41 05 23.78 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
