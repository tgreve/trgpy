
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-04-05T06:25:50PDT



Photometric Data for MM J18423+5938

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|MIPS 24 microns     |     |<0.6    |mJy                 |1.25E+13|        |0.6E-03|Jy|1990IRASF.C...0000M|3sigma uncertainty| 25        microns   | Broad-band measurement|115813.1 +302058 (B1950)| Flux in fixed aperture|                                        |From new raw data
2|IRAS 60 microns     |     |<100.   |mJy                 |5.00E+12|        |100.E-03|Jy|1990IRASF.C...0000M|3sigma uncertainty| 60        microns   | Broad-band measurement|115813.1 +302058 (B1950)| Flux in fixed aperture|IRAS quality flag = 3                   |From new raw data
3|MIPS 70 microns     | 31. | 4.     |mJy                 |4.28E+12|31.E-03 |+/-4.E-03|Jy|1990IRASF.C...0000M|uncertainty| 60        microns   | Broad-band measurement|115813.1 +302058 (B1950)| Flux in fixed aperture|IRAS quality flag = 3                   |From new raw data
4|IRAS 100 microns    |     |<6000.  |mJy                 |3.00E+12|        |600.E-03|Jy|1990IRASF.C...0000M|3sigma uncertainty| 100       microns   | Broad-band measurement|115813.1 +302058 (B1950)| Flux in fixed aperture|IRAS quality flag = 2                   |From new raw data
8|1.2 mm (MAMBO)      | 30  |+/-2    |milliJy             |2.50E+11|  3.00E-02|+/-2.00E-03|Jy|2010A&A...522L...4L|uncertainty|       1.2 mm        | Broad-band measurement|18 42 22.5 +59 38 30 (J2000)| Flux integrated from map|                                        |From new raw data
9|2 mm (EMIR)         | 9   |+/-3    |milliJy             |1.50E+11|  9.00E-03|+/-3.00E-03|Jy|2010A&A...522L...4L|uncertainty|         2 mm        | Broad-band measurement|18 42 22.5 +59 38 30 (J2000)| Flux integrated from map|                                        |From new raw data
10|3 mm (EMIR)        | 2   |+/-1.5  |milliJy             |0.99E+11|  2.00E-03|+/-1.50E-03|Jy|2010A&A...522L...4L|uncertainty|         3 mm        | Broad-band measurement|18 42 22.5 +59 38 30 (J2000)| Flux integrated from map|                                        |From new raw data
11|1.4GHz (VLA)       |     |<2.5    |milliJy             |1.40E+09|        |2.5E-03 |Jy|1995ApJ...450..559B|1sigma uncertainty reported|1.4        GHz       | Broad-band measurement; synthetic band|120046.812 +300414.82 (J2000)| From fitting to map|                                        |From new raw data; Corrected for contaminating sources
