
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-03-28T04:01:20PDT



Photometric Data for SMMJ02396-0134

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|3.6 microns (IRAC)  | 6.0704E+02|+/-1.0926E-01|microJy             |8.44E+13|  6.07E-04|+/-1.09E-07|Jy|2013SSTSLC4.2....0C|uncertainty|3.55       microns   | Broad-band measurement|| Flux in fixed aperture|5.8" aperture                           |From new raw data
4|4.5 microns (IRAC)  | 5.8006E+02|+/-1.0911E-01|microJy             |6.67E+13|  5.80E-04|+/-1.09E-07|Jy|2013SSTSLC4.2....0C|uncertainty|4.493      microns   | Broad-band measurement|| Flux in fixed aperture|5.8" aperture                           |From new raw data
5|5.8 microns (IRAC)  | 4.8860E+02|+/-4.2388E-01|microJy             |5.23E+13|  4.89E-04|+/-4.24E-07|Jy|2013SSTSLC4.2....0C|uncertainty|5.731      microns   | Broad-band measurement|| Flux in fixed aperture|5.8" aperture                           |From new raw data
8|8.0 microns (IRAC)  | 5.7169E+02|+/-7.3744E-01|microJy             |3.81E+13|  5.72E-04|+/-7.37E-07|Jy|2013SSTSLC4.2....0C|uncertainty|7.872      microns   | Broad-band measurement|| Flux in fixed aperture|5.8" aperture                           |From new raw data
9|24 microns (MIPS)   | 2.5121E+03|+/-1.9017E+01|microJy             |1.27E+13|  2.51E-03|+/-1.90E-05|Jy|2013SSTSLC4.2....0C|uncertainty|23.68      microns   | Broad-band measurement|| Modelled datum|PSF fit                                 |From new raw data
10|24 microns (MIPS)   | 2.4807E+03|+/-1.7395E+01|microJy             |1.27E+13|  2.48E-03|+/-1.74E-05|Jy|2013SSTSLC4.2....0C|uncertainty|23.68      microns   | Broad-band measurement|| Flux in fixed aperture|14.7" aperture                          |From new raw data
5|350 microns (SHARC2)| 51.0      |+/-6.0  |milliJy             |8.57E+11|  51.0E-03|+/-6.0E-03|Jy|2006ApJ...650..592K|uncertainty|     350   microns   | Broad-band measurement| | Total flux|                                        |From new raw data
6|450 microns (SCUBA) | 42.0      |+/-10   |milliJy             |6.66E+11|  42.0E-03|+/-10.0E-03|Jy|2007MNRAS.376.1073Z|uncertainty|     450   microns   | Broad-band measurement|02 39 56.3 -01 34 25 (J2000)| Flux integrated from map|                                        |From reprocessed raw data
6|450 microns (SCUBA) | 1.0       |+/-12   |milliJy             |6.66E+11|  1.0E-03|+/-12.0E-03|Jy|2007MNRAS.376.1073Z|uncertainty|     450   microns   | Broad-band measurement|02 39 56.3 -01 34 25 (J2000)| Flux integrated from map|                                        |From reprocessed raw data
11|450 microns (SCUBA) | 6         |+/-6    |milliJy             |6.66E+11|  6.00E-03|+/-6.00E-03|Jy|2007MNRAS.376.1073Z|uncertainty|     450   microns   | Broad-band measurement|02 39 56.3 -01 34 25 (J2000)| Flux integrated from map|                                        |From reprocessed raw data
7|850 microns (SCUBA) | 11.0      |+/-1.9  |milliJy             |3.53E+11|  11.0E-03|+/-1.9E-03|Jy|2007MNRAS.376.1073Z|uncertainty|     850   microns   | Broad-band measurement|02 39 56.3 -01 34 25 (J2000)| Flux integrated from map|S/N = 6.5                               |From reprocessed raw data
7|850 microns (SCUBA) | 6.8       |+/-0.9  |milliJy             |3.53E+11|  6.8E-03|+/-0.9E-03|Jy|2007MNRAS.376.1073Z|uncertainty|     850   microns   | Broad-band measurement|02 39 56.3 -01 34 25 (J2000)| Flux integrated from map|S/N = 6.5                               |From reprocessed raw data
7|850 microns (SCUBA) | 6.68      |+/-0.58 |milliJy             |3.53E+11|  6.68E-03|+/-0.58E-03|Jy|2007MNRAS.376.1073Z|uncertainty|     850   microns   | Broad-band measurement|02 39 56.3 -01 34 25 (J2000)| Flux integrated from map|S/N = 6.5                               |From reprocessed raw data
12|850 microns (SCUBA) | 6.2       ||milliJy             |3.53E+11|  6.20E-03||Jy|2007MNRAS.376.1073Z|no uncertainty reported|     850   microns   | Broad-band measurement|02 39 56.3 -01 34 25 (J2000)| Flux integrated from map|S/N = 6.5                               |From reprocessed raw data
7|880 microns (SMA)   | 7.95      |+/-0.60 |milliJy             |3.40E+11|  7.95E-03|+/-0.60E-03|Jy|2007MNRAS.376.1073Z|uncertainty|     850   microns   | Broad-band measurement|02 39 56.3 -01 34 25 (J2000)| Flux integrated from map|S/N = 6.5                               |From reprocessed raw data
27|1.4 GHz (VLA)      | 573.      |+/-11   |microJy             |1.40E+09|  573.E-06|+/-1.10E-05|Jy|2006MNRAS.371..963B|1 sigma|       1.4 GHz       | Broad-band measurement|16 36 58.179 +41 05 23.78 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
