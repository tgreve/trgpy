
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-07-10T08:18:23PDT



Photometric Data for SHADES J021738-050523

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|B (Subaru) AB       | 25.36     |+/-0.01 |mag                 |6.69E+14|  2.61E-07|+/-2.40E-09|Jy|2008MNRAS.387..247C|uncertainty|      4478 A         | Broad-band measurement|34.412021 -5.091103 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
2|V (Subaru) AB       | 24.85     |+/-0.01 |mag                 |5.46E+14|  4.17E-07|+/-3.84E-09|Jy|2008MNRAS.387..247C|uncertainty|      5493 A         | Broad-band measurement|34.412021 -5.091103 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
3|R (Subaru) AB       | 24.59     |+/-0.01 |mag                 |4.58E+14|  5.30E-07|+/-4.88E-09|Jy|2008MNRAS.387..247C|uncertainty|      6550 A         | Broad-band measurement|34.412021 -5.091103 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
4|i' (Subaru) AB      | 24.39     |+/-0.01 |mag                 |3.89E+14|  6.37E-07|+/-5.86E-09|Jy|2008MNRAS.387..247C|uncertainty|      7709 A         | Broad-band measurement|34.412021 -5.091103 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
5|z' (Subaru) AB      | 24.05     |+/-0.02 |mag                 |3.31E+14|  8.71E-07|+/-1.60E-08|Jy|2008MNRAS.387..247C|uncertainty|      9054 A         | Broad-band measurement|34.412021 -5.091103 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
6|3.6 microns (IRAC)  | 2.2515E+01|+/-1.0165E-01|microJy             |8.44E+13|  2.25E-05|+/-1.02E-07|Jy|2013SSTSLC4.2....0C|uncertainty|3.55       microns   | Broad-band measurement|| Flux in fixed aperture|3.8" aperture                           |From new raw data
7|3.6 microns (IRAC)  | 2.4189E+01|+/-6.3391E-01|microJy             |8.44E+13|  2.42E-05|+/-6.34E-07|Jy|2013SSTSLC4.2....0C|uncertainty|3.55       microns   | Broad-band measurement|| Flux in fixed aperture|3.8" aperture                           |From new raw data
8|3.6 microns (IRAC)  | 3.0532E+01|+/-1.3104E-01|microJy             |8.44E+13|  3.05E-05|+/-1.31E-07|Jy|2013SSTSLC4.2....0C|uncertainty|3.55       microns   | Broad-band measurement|| Flux in fixed aperture|5.8" aperture                           |From new raw data
9|3.6 microns (IRAC)  | 3.4384E+01|+/-1.0264E+00|microJy             |8.44E+13|  3.44E-05|+/-1.03E-06|Jy|2013SSTSLC4.2....0C|uncertainty|3.55       microns   | Broad-band measurement|| Flux in fixed aperture|5.8" aperture                           |From new raw data
6|3.6 microns (IRAC)  | 25.19     |+/-0.85 | microJy            |8.44E+13|  2.52E-05|+/-8.50E-07|Jy|2008MNRAS.387..247C|uncertainty|     3.550 microns   | Broad-band measurement|34.412021 -5.091103 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
11|4.5 microns (IRAC)  | 3.7630E+01|+/-2.6744E-01|microJy             |6.67E+13|  3.76E-05|+/-2.67E-07|Jy|2013SSTSLC4.2....0C|uncertainty|4.493      microns   | Broad-band measurement|| Flux in fixed aperture|5.8" aperture                           |From new raw data
12|4.5 microns (IRAC)  | 3.6014E+01|+/-1.7305E+00|microJy             |6.67E+13|  3.60E-05|+/-1.73E-06|Jy|2013SSTSLC4.2....0C|uncertainty|4.493      microns   | Broad-band measurement|| Flux in fixed aperture|5.8" aperture                           |From new raw data
13|4.5 microns (IRAC)  | 2.7662E+01|+/-1.0689E+00|microJy             |6.67E+13|  2.77E-05|+/-1.07E-06|Jy|2013SSTSLC4.2....0C|uncertainty|4.493      microns   | Broad-band measurement|| Flux in fixed aperture|3.8" aperture                           |From new raw data
14|4.5 microns (IRAC)  | 2.8849E+01|+/-1.8128E-01|microJy             |6.67E+13|  2.88E-05|+/-1.81E-07|Jy|2013SSTSLC4.2....0C|uncertainty|4.493      microns   | Broad-band measurement|| Flux in fixed aperture|3.8" aperture                           |From new raw data
7|4.5 microns (IRAC)  | 29.02     |+/-1.19 | microJy            |6.67E+13|  2.90E-05|+/-1.19E-06|Jy|2008MNRAS.387..247C|uncertainty|     4.493 microns   | Broad-band measurement|34.412021 -5.091103 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
16|5.8 microns (IRAC)  | 5.1453E+01|+/-4.1953E+00|microJy             |5.23E+13|  5.15E-05|+/-4.20E-06|Jy|2013SSTSLC4.2....0C|uncertainty|5.731      microns   | Broad-band measurement|| Flux in fixed aperture|3.8" aperture                           |From new raw data
17|5.8 microns (IRAC)  | 7.0967E+01|+/-6.3387E+00|microJy             |5.23E+13|  7.10E-05|+/-6.34E-06|Jy|2013SSTSLC4.2....0C|uncertainty|5.731      microns   | Broad-band measurement|| Flux in fixed aperture|5.8" aperture                           |From new raw data
18|5.8 microns (IRAC)  | 4.1171E+01|+/-4.9339E-01|microJy             |5.23E+13|  4.12E-05|+/-4.93E-07|Jy|2013SSTSLC4.2....0C|uncertainty|5.731      microns   | Broad-band measurement|| Flux in fixed aperture|3.8" aperture                           |From new raw data
19|5.8 microns (IRAC)  | 5.0153E+01|+/-6.4457E-01|microJy             |5.23E+13|  5.02E-05|+/-6.45E-07|Jy|2013SSTSLC4.2....0C|uncertainty|5.731      microns   | Broad-band measurement|| Flux in fixed aperture|5.8" aperture                           |From new raw data
8|5.8 microns (IRAC)  | 47.81     |+/-5.50 | microJy            |5.23E+13|  4.78E-05|+/-5.50E-06|Jy|2008MNRAS.387..247C|uncertainty|     5.731 microns   | Broad-band measurement|34.412021 -5.091103 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
9|15 microns (AKARI)  | 35        |+/-19   |microJy             |1.92E+13|  3.50E-05|+/-1.90E-05|Jy|2010A&A...514A..10S|uncertainty|     15.58 microns   | Broad-band measurement|| Flux in fixed aperture|                                        |From new raw data
10|24 microns (MIPS)   | 325.0     |+/-47.0 | microJy            |1.27E+13|  3.25E-04|+/-4.70E-05|Jy|2007MNRAS.380..199I|rms uncertainty|     23.68 microns   | Broad-band measurement|02 17 38.86 -05 05 29.1 (J2000)| Flux integrated from map|                                        |Averaged from previously published data
11|24 microns (MIPS)   | 303.42    |+/-18.84| microJy            |1.27E+13|  3.03E-04|+/-1.88E-05|Jy|2008MNRAS.387..247C|uncertainty|     23.68 microns   | Broad-band measurement|34.412021 -5.091103 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
28|24 microns (MIPS)   | 3.5048E+02|+/-1.2341E+01|microJy             |1.27E+13|  3.50E-04|+/-1.23E-05|Jy|2013SSTSLC4.2....0C|uncertainty|23.68      microns   | Broad-band measurement|| Modelled datum|PSF fit                                 |From new raw data
29|24 microns (MIPS)   | 3.0441E+02|+/-6.0882E+01|microJy             |1.27E+13|  3.04E-04|+/-6.09E-05|Jy|2013SSTSLC4.2....0C|uncertainty|23.68      microns   | Broad-band measurement|| Modelled datum|PSF fit                                 |From new raw data
30|24 microns (MIPS)   | 3.9182E+02|+/-1.1789E+01|microJy             |1.27E+13|  3.92E-04|+/-1.18E-05|Jy|2013SSTSLC4.2....0C|uncertainty|23.68      microns   | Broad-band measurement|| Flux in fixed aperture|14.7" aperture                          |From new raw data
31|24 microns (MIPS)   | 3.2324E+02|+/-5.7965E+01|microJy             |1.27E+13|  3.23E-04|+/-5.80E-05|Jy|2013SSTSLC4.2....0C|uncertainty|23.68      microns   | Broad-band measurement|| Flux in fixed aperture|14.7" aperture                          |From new raw data
1|250 microns (SPIRE) | 24.8     |+/-3.6  |mJy |1.199e+12|24.8E-03  |+/-3.6E-03  |Jy|Reference          |uncertainty       | | | | |
2|350 microns (SPIRE) | 26.2     |+/-4.2  |mJy |8.57e+11|26.2E-03   |+/-4.2E-03  |Jy|Reference          |uncertainty       | | | | |
3|500 microns (SPIRE) | 26.0     |+/-4.8  |mJy |5.996e+11|26.0E-03  |+/-4.8E-03  |Jy|Reference          |uncertainty       | | | | |
12|850 microns (SCUBA) | 7.1       |+/-1.5  | milliJy            |3.53E+11|  7.10E-03|+/-1.50E-03|Jy|2008MNRAS.387..247C|uncertainty|       850 microns   | Broad-band measurement|34.412021 -5.091103 (J2000)| Flux integrated from map|                                        |Averaged from previously published data
13|850 microns (SCUBA) | 7.1       |+/-1.6  | milliJy            |3.53E+11|  7.10E-03|+/-1.60E-03|Jy|2007MNRAS.380..199I|rms uncertainty|       850 microns   | Broad-band measurement|02 17 38.921 -05 05 23.72 (J2000)| Flux integrated from map|                                        |Averaged from previously published data
5|2.0 mm (PdBI)       | 0.3      |+/-0.1  |mJy |1.54E+11|0.3E-03|+/-0.1E-03|Jy|2010Natur.464..733S|uncertainty|       2.8 microns   | Broad-band measurement|21 35 11.6 -01 02 52.0 (J2000)| Flux in fixed aperture|                                        |From new raw data
6|1.4 GHz (VLA)       | 57       |+/-10   |uJy |1.40E+09|57.E-06|+/-10.E-06|Jy|2006MNRAS.371..963B|1 sigma|       1.4 GHz       | Broad-band measurement|16 36 55.767 +40 59 09.97 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
14|1.4 GHz (VLA)       | 41.2      |+/-11.3 |microJy             |1.40E+09|  4.12E-05|+/-1.13E-05|Jy|2007MNRAS.380..199I|rms uncertainty|       1.4 GHz       | Broad-band measurement|02 17 38.878 -05 05 28.03 (J2000)| Flux integrated from map|                                        |From new raw data
