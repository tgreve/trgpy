
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-07-10T04:03:58PDT



Photometric Data for 2MASSi J1005174+434609

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|FUV (GALEX) AB      | 19.047    |+/-0.116|mag                 |1.97E+15|  8.73E-05|+/-9.33E-06|Jy|2007AJ....133.1780T|uncertainty|    1525   A         | Broad-band measurement|151.322624 43.769218 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
2|FUV (GALEX) AB      | 19.1973   |+/-0.136245|mag                 |1.95E+15|  7.61E-05|+/-9.54E-06|Jy|2012GASC..C...0000S|uncertainty|1538.6     A         | Broad-band measurement|151.32264688452 43.769284024179 (J2000)| Flux integrated from map|Kron flux in elliptical aperture        |From new raw data
3|FUV (GALEX) AB      | 19.4514   |+/-0.159697|mag                 |1.95E+15|  6.02E-05|+/-8.85E-06|Jy|2012GASC..C...0000S|uncertainty|1538.6     A         | Broad-band measurement|151.32264688452 43.769284024179 (J2000)| Flux in fixed aperture|Flux in 7.5 arcsec diameter aperture    |From new raw data
4|1700 A (SDSS)       | -14.588   ||log(erg/cm^2^/s/A)  |1.76E+15|  2.49E-04||Jy|2011MNRAS.410..860A|no uncertainty reported|      1700 A         | Broad-band measurement|151.322632 +43.769253 (J2000)| Flux integrated from map|                                        |From reprocessed raw data
5|NUV (GALEX) AB      | 18.387    |+/-0.048|mag                 |1.36E+15|  1.60E-04|+/-7.09E-06|Jy|2007AJ....133.1780T|uncertainty|    2200   A         | Broad-band measurement|151.322624 43.769218 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
6|NUV (GALEX) AB      | 18.4957   |+/-0.0572784|mag                 |1.29E+15|  1.45E-04|+/-7.65E-06|Jy|2012GASC..C...0000S|uncertainty|2315.7     A         | Broad-band measurement|151.32264688452 43.769284024179 (J2000)| Flux integrated from map|Kron flux in elliptical aperture        |From new raw data
7|NUV (GALEX) AB      | 18.9286   |+/-0.0749882|mag                 |1.29E+15|  9.74E-05|+/-6.73E-06|Jy|2012GASC..C...0000S|uncertainty|2315.7     A         | Broad-band measurement|151.32264688452 43.769284024179 (J2000)| Flux in fixed aperture|Flux in 7.5 arcsec diameter aperture    |From new raw data
8|u (SDSS CModel) AB  | 16.986    ||asinh mag           |8.36E+14|  5.83E-04||Jy|2004SDSS3.C...0000:|no uncertainty reported|3585       A         | Broad-band measurement|151.322632 43.769249 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; PETROFAINT - Petrosian radius measured at very low surface brightness; TOO_LARGE - very large object, poorly determined sky, or bad deblend; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
9|u (SDSS Petrosian)AB| 17.040    |+/-0.007|asinh mag           |8.36E+14|  5.76E-04|+/-3.59E-06|Jy|2004SDSS3.C...0000:|based on count statistics only|3585       A         | Broad-band measurement|151.322632 43.769249 (J2000)| Modelled datum|From new raw data
10|u (SDSS PSF) AB     | 16.980    |+/-0.021|asinh mag           |8.36E+14|  6.08E-04|+/-1.16E-05|Jy|2004SDSS3.C...0000:|based on count statistics only|3585       A         | Broad-band measurement|151.322632 43.769249 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; PETROFAINT - Petrosian radius measured at very low surface brightness; TOO_LARGE - very large object, poorly determined sky, or bad deblend; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
11|u (SDSS PSF) AB     | 16.980    |+/-0.021|asinh mag           |8.36E+14|  6.08E-04|+/-1.18E-05|Jy|2007SDSS6.C...0000:|based on count statistics only|3585       A         | Broad-band measurement|151.3226311778 43.7692517886 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; PETROFAINT - Petrosian radius measured at very low surface brightness; TOO_LARGE - very large object, poorly determined sky, or bad deblend; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
12|u (SDSS Model) AB   | 16.985    |+/-0.007|asinh mag           |8.36E+14|  6.05E-04|+/-4.14E-06|Jy|2004SDSS3.C...0000:|based on count statistics only|3585       A         | Broad-band measurement|151.322632 43.769249 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; PETROFAINT - Petrosian radius measured at very low surface brightness; TOO_LARGE - very large object, poorly determined sky, or bad deblend; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
13|g (SDSS Petrosian)AB| 16.851    |+/-0.003|asinh mag           |6.17E+14|  6.60E-04|+/-1.78E-06|Jy|2004SDSS3.C...0000:|based on count statistics only|4858       A         | Broad-band measurement|151.322632 43.769249 (J2000)| Modelled datum|From new raw data
14|g (SDSS PSF) AB     | 16.776    |+/-0.031|asinh mag           |6.17E+14|  7.07E-04|+/-2.02E-05|Jy|2007SDSS6.C...0000:|based on count statistics only|4858       A         | Broad-band measurement|151.3226311778 43.7692517886 (J2000)| Modelled datum|SDSS flags: MANYPETRO - more than one Petrosian radius; BAD_RADIAL - some low S/N radial points; TOO_LARGE - very large object, poorly determined sky, or bad deblend; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
15|g (SDSS CModel) AB  | 16.803    ||asinh mag           |6.17E+14|  6.90E-04||Jy|2004SDSS3.C...0000:|no uncertainty reported|4858       A         | Broad-band measurement|151.322632 43.769249 (J2000)| Modelled datum|SDSS flags: MANYPETRO - more than one Petrosian radius; BAD_RADIAL - some low S/N radial points; TOO_LARGE - very large object, poorly determined sky, or bad deblend; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
16|g (SDSS PSF) AB     | 16.776    |+/-0.031|asinh mag           |6.17E+14|  7.08E-04|+/-2.02E-05|Jy|2004SDSS3.C...0000:|based on count statistics only|4858       A         | Broad-band measurement|151.322632 43.769249 (J2000)| Modelled datum|SDSS flags: MANYPETRO - more than one Petrosian radius; BAD_RADIAL - some low S/N radial points; TOO_LARGE - very large object, poorly determined sky, or bad deblend; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
17|g (SDSS Model) AB   | 16.803    |+/-0.004|asinh mag           |6.17E+14|  6.90E-04|+/-2.67E-06|Jy|2004SDSS3.C...0000:|based on count statistics only|4858       A         | Broad-band measurement|151.322632 43.769249 (J2000)| Modelled datum|SDSS flags: MANYPETRO - more than one Petrosian radius; BAD_RADIAL - some low S/N radial points; TOO_LARGE - very large object, poorly determined sky, or bad deblend; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
18|r (SDSS CModel) AB  | 16.631    ||asinh mag           |4.77E+14|  8.09E-04||Jy|2004SDSS3.C...0000:|no uncertainty reported|6290       A         | Broad-band measurement|151.322632 43.769249 (J2000)| Modelled datum|SDSS flags: MANYPETRO - more than one Petrosian radius; BAD_RADIAL - some low S/N radial points; TOO_LARGE - very large object, poorly determined sky, or bad deblend; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding; CANONICAL_BAND - this band was primary (usually r);|From new raw data
19|r (SDSS Petrosian)AB| 16.680    |+/-0.003|asinh mag           |4.77E+14|  7.72E-04|+/-2.03E-06|Jy|2004SDSS3.C...0000:|based on count statistics only|6290       A         | Broad-band measurement|151.322632 43.769249 (J2000)| Modelled datum|From new raw data
20|r (SDSS Model) AB   | 16.631    |+/-0.004|asinh mag           |4.77E+14|  8.09E-04|+/-3.21E-06|Jy|2004SDSS3.C...0000:|based on count statistics only|6290       A         | Broad-band measurement|151.322632 43.769249 (J2000)| Modelled datum|SDSS Effective Radius =   0.02" x   0.01".;SDSS flags: MANYPETRO - more than one Petrosian radius; BAD_RADIAL - some low S/N radial points; TOO_LARGE - very large object, poorly determined sky, or bad deblend; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding; CANONICAL_BAND - this band was primary (usually r);|From new raw data
21|r (SDSS PSF) AB     | 16.637    |+/-0.017|asinh mag           |4.77E+14|  8.04E-04|+/-1.26E-05|Jy|2007SDSS6.C...0000:|based on count statistics only|6290       A         | Broad-band measurement|151.3226311778 43.7692517886 (J2000)| Modelled datum|SDSS flags: MANYPETRO - more than one Petrosian radius; BAD_RADIAL - some low S/N radial points; TOO_LARGE - very large object, poorly determined sky, or bad deblend; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding; CANONICAL_BAND - this band was primary (usually r);|From new raw data
22|r (SDSS PSF) AB     | 16.637    |+/-0.017|asinh mag           |4.77E+14|  8.04E-04|+/-1.26E-05|Jy|2004SDSS3.C...0000:|based on count statistics only|6290       A         | Broad-band measurement|151.322632 43.769249 (J2000)| Modelled datum|SDSS flags: MANYPETRO - more than one Petrosian radius; BAD_RADIAL - some low S/N radial points; TOO_LARGE - very large object, poorly determined sky, or bad deblend; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding; CANONICAL_BAND - this band was primary (usually r);|From new raw data
23|i (SDSS Petrosian)AB| 16.522    |+/-0.003|asinh mag           |3.89E+14|  1.45E-03|+/-4.43E-06|Jy|2004SDSS3.C...0000:|based on count statistics only|7706       A         | Broad-band measurement|151.322632 43.769249 (J2000)| Modelled datum|From new raw data
24|i (SDSS CModel) AB  | 16.469    ||asinh mag           |3.89E+14|  9.38E-04||Jy|2004SDSS3.C...0000:|no uncertainty reported|7706       A         | Broad-band measurement|151.322632 43.769249 (J2000)| Modelled datum|SDSS flags: MANYPETRO - more than one Petrosian radius; BAD_RADIAL - some low S/N radial points; TOO_LARGE - very large object, poorly determined sky, or bad deblend; ELLIPFAINT - no isophotal fits performed; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
25|i (SDSS PSF) AB     | 16.482    |+/-0.015|asinh mag           |3.89E+14|  9.27E-04|+/-1.28E-05|Jy|2007SDSS6.C...0000:|based on count statistics only|7706       A         | Broad-band measurement|151.3226311778 43.7692517886 (J2000)| Modelled datum|SDSS flags: MANYPETRO - more than one Petrosian radius; BAD_RADIAL - some low S/N radial points; TOO_LARGE - very large object, poorly determined sky, or bad deblend; ELLIPFAINT - no isophotal fits performed; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
26|i (SDSS PSF) AB     | 16.482    |+/-0.015|asinh mag           |3.89E+14|  9.28E-04|+/-1.32E-05|Jy|2004SDSS3.C...0000:|based on count statistics only|7706       A         | Broad-band measurement|151.322632 43.769249 (J2000)| Modelled datum|SDSS flags: MANYPETRO - more than one Petrosian radius; BAD_RADIAL - some low S/N radial points; TOO_LARGE - very large object, poorly determined sky, or bad deblend; ELLIPFAINT - no isophotal fits performed; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
27|i (SDSS Model) AB   | 16.469    |+/-0.005|asinh mag           |3.89E+14|  9.39E-04|+/-3.96E-06|Jy|2004SDSS3.C...0000:|based on count statistics only|7706       A         | Broad-band measurement|151.322632 43.769249 (J2000)| Modelled datum|SDSS flags: MANYPETRO - more than one Petrosian radius; BAD_RADIAL - some low S/N radial points; TOO_LARGE - very large object, poorly determined sky, or bad deblend; ELLIPFAINT - no isophotal fits performed; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
28|z (SDSS PSF) AB     | 16.251    |+/-0.020|asinh mag           |3.25E+14|  1.13E-03|+/-2.07E-05|Jy|2007SDSS6.C...0000:|based on count statistics only|9222       A         | Broad-band measurement|151.3226311778 43.7692517886 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; TOO_LARGE - very large object, poorly determined sky, or bad deblend; ELLIPFAINT - no isophotal fits performed; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
29|z (SDSS Petrosian)AB| 16.292    |+/-0.008|asinh mag           |3.25E+14|  1.08E-03|+/-7.76E-06|Jy|2004SDSS3.C...0000:|based on count statistics only|9222       A         | Broad-band measurement|151.322632 43.769249 (J2000)| Modelled datum|From new raw data
30|z (SDSS CModel) AB  | 16.250    ||asinh mag           |3.25E+14|  1.15E-03||Jy|2004SDSS3.C...0000:|no uncertainty reported|9222       A         | Broad-band measurement|151.322632 43.769249 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; TOO_LARGE - very large object, poorly determined sky, or bad deblend; ELLIPFAINT - no isophotal fits performed; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
31|z (SDSS PSF) AB     | 16.251    |+/-0.020|asinh mag           |3.25E+14|  1.13E-03|+/-2.04E-05|Jy|2004SDSS3.C...0000:|based on count statistics only|9222       A         | Broad-band measurement|151.322632 43.769249 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; TOO_LARGE - very large object, poorly determined sky, or bad deblend; ELLIPFAINT - no isophotal fits performed; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
32|z (SDSS Model) AB   | 16.249    |+/-0.007|asinh mag           |3.25E+14|  1.13E-03|+/-7.49E-06|Jy|2004SDSS3.C...0000:|based on count statistics only|9222       A         | Broad-band measurement|151.322632 43.769249 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; TOO_LARGE - very large object, poorly determined sky, or bad deblend; ELLIPFAINT - no isophotal fits performed; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
33|J (2MASS)           | 1.02e-03  || Jy                 |2.40E+14|  1.02E-03||Jy|2008MNRAS.383.1513L|no uncertainty reported|      1.25 microns   | Broad-band measurement|10 05 17.43 +43 46 09.3 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data; Extinction-correctedfor Milky Way
34|H (2MASS)           | 9.73e-04  || Jy                 |1.82E+14|  9.73E-04||Jy|2008MNRAS.383.1513L|no uncertainty reported|      1.65 microns   | Broad-band measurement|10 05 17.43 +43 46 09.3 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data; Extinction-correctedfor Milky Way
35|K_s (2MASS)         | 1.30e-03  || Jy                 |1.38E+14|  1.30E-03||Jy|2008MNRAS.383.1513L|no uncertainty reported|      2.17 microns   | Broad-band measurement|10 05 17.43 +43 46 09.3 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data; Extinction-correctedfor Milky Way
36|350 microns SHARC II| 77        |+/-14   |milliJy             |8.57E+11|  7.70E-02|+/-1.40E-02|Jy|2006ApJ...642..694B|1 sigma|     350   microns   | Broad-band measurement|10 05 17.45 +43 46 09.30 (J2000)| Flux integrated from map|                                        |From new raw data
37|1.2 mm (MAMBO)      | 4.2       |+/-0.8  | milliJy            |2.50E+11|  4.20E-03|+/-8.00E-04|Jy|2003A&A...398..857O|uncertainty|       1.2 mm        | Broad-band measurement|10 05 17.5 +43 46 09.0 (J2000)| Flux integrated from map|                                        |From new raw data
