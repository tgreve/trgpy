
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-06-16T16:23:52PDT



Photometric Data for DEEP2 13017843

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|5-10 keV (Chandra)  ||<0.60E-15  |erg/cm^2^/s         |1.81E+18||3.31E-11|Jy|2009ApJS..180..102L|1 sigma|      7.50 keV       | Broad-band measurement|215.079029 +52.934240 (J2000)| Modelled datum|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
2|2-10 keV (Chandra)  ||<0.49E-15  |erg/cm^2^/s         |1.45E+18||3.38E-11|Jy|2009ApJS..180..102L|1 sigma|      6.00 keV       | Broad-band measurement|215.079029 +52.934240 (J2000)| Modelled datum|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
3|0.5-10 keV (Chandra)| 0.98E-15  |+/-0.44E-15|erg/cm^2^/s         |1.27E+18|  7.72E-11|+/-3.46E-11|Jy|2009ApJS..180..102L|1 sigma|      5.25 keV       | Broad-band measurement|215.079029 +52.934240 (J2000)| Modelled datum|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
4|0.5-2 keV (Chandra) | 0.48E-15  |+/-0.14E-15|erg/cm^2^/s         |3.02E+17|  1.59E-10|+/-4.64E-11|Jy|2009ApJS..180..102L|1 sigma|      1.25 keV       | Broad-band measurement|215.079029 +52.934240 (J2000)| Modelled datum|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
5|K_s (Keck)          | 18.67     || mag                |1.39E+14|  2.11E-05||Jy|2007MNRAS.382..109T|no uncertainty reported|      2.15 microns   | Broad-band measurement|215.07828 +52.93483 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
