
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-06-17T08:38:21PDT



Photometric Data for IOK 1

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
3|i' (Subaru) AB      ||>27.84     |mag                 |3.89E+14||2.66E-08|Jy|2008ApJ...677...12O|2 sigma|      7709 A         | Broad-band measurement|13 23 59.8 +27 24 55.8 (J2000)| Flux in fixed aperture|2" aperture                             |From reprocessed raw data
4|NB816 (Subaru) AB   ||>27.04     |mag                 |3.68E+14||5.55E-08|Jy|2008ApJ...677...12O|2 sigma|      8150 A         | Broad-band measurement|13 23 59.8 +27 24 55.8 (J2000)| Flux in fixed aperture|2" aperture                             |From reprocessed raw data
5|z' (Subaru) AB      ||>27.04     |mag                 |3.31E+14||5.55E-08|Jy|2008ApJ...677...12O|2 sigma|      9054 A         | Broad-band measurement|13 23 59.8 +27 24 55.8 (J2000)| Flux in fixed aperture|2" aperture                             |From reprocessed raw data
6|NB921 (Subaru) AB   ||>26.96     |mag                 |3.26E+14||5.97E-08|Jy|2008ApJ...677...12O|2 sigma|      9196 A         | Broad-band measurement|13 23 59.8 +27 24 55.8 (J2000)| Flux in fixed aperture|2" aperture                             |From reprocessed raw data
7|NB973 (Subaru) AB   | 24.40     ||mag                 |3.07E+14|  6.31E-07||Jy|2008ApJ...677...12O|no uncertainty reported|      9755 A         | Broad-band measurement|13 23 59.8 +27 24 55.8 (J2000)| Total flux|                                        |From new raw data
8|NB973 (Subaru) AB   | 24.60     ||mag                 |3.07E+14|  5.25E-07||Jy|2008ApJ...677...12O|no uncertainty reported|      9755 A         | Broad-band measurement|13 23 59.8 +27 24 55.8 (J2000)| Flux in fixed aperture|2" aperture                             |From new raw data
9|y (Subaru) AB       | 25.42     ||mag                 |3.04E+14|  2.47E-07||Jy|2009ApJ...706.1136O|no uncertainty reported|      9860 A         | Broad-band measurement|| Flux in fixed aperture|1.8" diameter aperture                  |From new raw data; Extinction-corrected for Milky Way
10|F125W (HST WFC3) AB      | 25.59     |+/-0.05 |mag                 |2.40E+14|  2.11E-07|+/-9.71E-09|Jy|2011ApJ...736L..28C|uncertainty|     12486 A         | Broad-band measurement|| Flux in fixed aperture|                                        |From new raw data
11|F130N (HST WFC3) AB      | 25.42     |+/-0.17 |mag                 |2.31E+14|  2.47E-07|+/-3.86E-08|Jy|2011ApJ...736L..28C|uncertainty|     13006 A         | Broad-band measurement|| Flux in fixed aperture|                                        |From new raw data
5|3.6 microns (IRAC)  |       |>23.99 |mag             |8.44E+13|  |9.205e-07|Jy|2010Natur.464..733S|3sigma uncertainty|     3.550 microns   | Broad-band measurement|21 35 11.6 -01 02 52.0 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
6|4.5 microns (IRAC)  |       |>23.54 |mag             |6.67E+13|  |1.393e-06|Jy|2010Natur.464..733S|3sigma uncertainty|     4.493 microns   | Broad-band measurement|21 35 11.6 -01 02 52.0 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
11|CARMA 238GHz      |      |<0.19 |mJy                 |2.39E+11|  |0.19E-03|Jy|2011ApJ...736L..28C|1sigma uncertainty|     13006 A         | Broad-band measurement|| Flux in fixed aperture|                                        |From new raw data
