
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-07-10T12:57:42PDT



Photometric Data for LEDA 2830631

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|Ly{alpha} (VLT)     | 2.9E-16   |+/-0.3E-16|erg s^-1^ cm^-2^    |2.47E+15|  2.90E+07|+/-3.00E+06|Jy-Hz|2007A&A...461..823V|uncertainty|    1216   A         | Line measurement; flux integrated over line; lines measured in emission|20 51 03.45 -27 03 04.1 (J2000)| From fitting to map|                                        |From new raw data
2|3.6 microns (IRAC)  | 59.5      |+/-6.2  | microJy            |8.44E+13|  5.95E-05|+/-6.20E-06|Jy|2007ApJS..171..353S|uncertainty|   3.550   microns   | Broad-band measurement|20 51 03.6 -27 03 02.53 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
3|4.5 microns (IRAC)  | 72.6      |+/-7.5  | microJy            |6.67E+13|  7.26E-05|+/-7.50E-06|Jy|2007ApJS..171..353S|uncertainty|   4.493   microns   | Broad-band measurement|20 51 03.6 -27 03 02.53 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
4|5.8 microns (IRAC)  | 78.3      |+/-10.4 | microJy            |5.23E+13|  7.83E-05|+/-1.04E-05|Jy|2007ApJS..171..353S|uncertainty|   5.731   microns   | Broad-band measurement|20 51 03.6 -27 03 02.53 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
5|8.0 microns (IRAC)  | 38.4      |+/-13.1 | microJy            |3.81E+13|  3.84E-05|+/-1.31E-05|Jy|2007ApJS..171..353S|uncertainty|   7.872   microns   | Broad-band measurement|20 51 03.6 -27 03 02.53 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
6|16 microns (IRS)    ||<141.0     | microJy            |1.87E+13||1.41E-04|Jy|2007ApJS..171..353S|3 sigma|      16   microns   | Broad-band measurement|20 51 03.6 -27 03 02.53 (J2000)| Flux in fixed aperture|6" diameter aperture                    |From reprocessed raw data
7|4.85 GHz            | 115       |+/-12   |milliJy             |4.85E+09|  1.15E-01|+/-1.20E-02|Jy|1994ApJS...90..179G|rms noise|4.85       GHz       | Broad-band measurement|205101.8 -270247 (J2000)| Modelled datum|                                        |From new raw data; Corrected for contaminating sources
8|1.4GHz (VLA)        | 498.1     |+/-15.0 |milliJy             |1.40E+09|  4.98E-01|+/-1.50E-02|Jy|1998AJ....115.1693C|uncertainty|    1.40   GHz       | Broad-band measurement|20 51 3.60 -27 03 3.1 (J2000)| Flux integrated from map|High peak                               |From new raw data
9|408 MHz             | 1.98      |+/-0.19 |Jy                  |4.08E+08|  1.98E+00|+/-1.90E-01|Jy|1981MNRAS.194..693L|rms noise|408        MHz       | Broad-band measurement|204805.0 -271426 (B1950)| Modelled datum|                                        |From new raw data; Corrected for contaminating sources
10|365 MHz (Texas)     | 2.255     |+/-0.056|Jy                  |3.65E+08|  2.25E+00|+/-5.60E-02|Jy|1996AJ....111.1945D|internal error|365        MHz       | Broad-band measurement; obtained by interpolation over frequency|204804.507 -271418.35 (B1950)| Integrated from scans|Model:P;MFlag:+;EFlag:+;LFlag:+.Poss var|From new raw data
