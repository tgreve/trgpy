
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-07-08T06:32:09PDT



Photometric Data for SDSS J123645.73+620754.4

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|4.0-8 keV (Chandra) ||<0.42E-15  |ergs cm^-2^ s^-1^   |1.45E+18||2.89E-11|Jy|2003AJ....126..539A|3 sigma|       6   keV       | Broad-band measurement|12 36 45.81 +62 07 53.9 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
2|4-8 keV (Chandra)   ||<0.57E-15  |erg cm^-2^ s^-1^    |1.45E+18||3.93E-11|Jy|2001AJ....122.2810B|no uncertainty reported|       6   keV       | Broad-band measurement|12 36 45.88 +62 07 54.1 (J2000)| Flux in fixed aperture|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
3|2-8 keV (Chandra)   ||<0.40E-15  |erg cm^-2^ s^-1^    |1.21E+18||3.31E-11|Jy|2001AJ....122.2810B|no uncertainty reported|       5   keV       | Broad-band measurement|12 36 45.88 +62 07 54.1 (J2000)| Flux in fixed aperture|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
4|2.0-8 keV (Chandra) ||<0.34E-15  |ergs cm^-2^ s^-1^   |1.21E+18||2.81E-11|Jy|2003AJ....126..539A|3 sigma|       5   keV       | Broad-band measurement|12 36 45.81 +62 07 53.9 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
5|0.5-8 keV (Chandra) | 0.20E-15  |+/-4   %|erg cm^-2^ s^-1^    |1.03E+18|  1.94E-11|+/-7.77E-13|Jy|2001AJ....122.2810B|estimated error|    4.25   keV       | Broad-band measurement|12 36 45.88 +62 07 54.1 (J2000)| Flux in fixed aperture|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
6|0.5-8 keV (Chandra) | 0.34E-15  ||ergs cm^-2^ s^-1^   |1.03E+18|  3.31E-11||Jy|2003AJ....126..539A|no uncertainty reported|    4.25   keV       | Broad-band measurement|12 36 45.81 +62 07 53.9 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
7|2.0-4 keV (Chandra) | 0.10E-15  ||ergs cm^-2^ s^-1^   |7.25E+17|  1.38E-11||Jy|2003AJ....126..539A|no uncertainty reported|       3   keV       | Broad-band measurement|12 36 45.81 +62 07 53.9 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
8|1.0-2 keV (Chandra) | 0.07E-15  ||ergs cm^-2^ s^-1^   |3.63E+17|  1.93E-11||Jy|2003AJ....126..539A|no uncertainty reported|     1.5   keV       | Broad-band measurement|12 36 45.81 +62 07 53.9 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
9|0.5-2 keV (Chandra) | 0.09E-15  ||ergs cm^-2^ s^-1^   |3.02E+17|  2.98E-11||Jy|2003AJ....126..539A|no uncertainty reported|    1.25   keV       | Broad-band measurement|12 36 45.81 +62 07 53.9 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
10|0.5-2 keV (Chandra) | 0.10E-15  |+/-4   %|erg cm^-2^ s^-1^    |3.02E+17|  3.31E-11|+/-1.32E-12|Jy|2001AJ....122.2810B|estimated error|    1.25   keV       | Broad-band measurement|12 36 45.88 +62 07 54.1 (J2000)| Flux in fixed aperture|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
11|0.5-1 keV (Chandra) ||<0.05E-15  |ergs cm^-2^ s^-1^   |1.81E+17||2.76E-11|Jy|2003AJ....126..539A|3 sigma|    0.75   keV       | Broad-band measurement|12 36 45.81 +62 07 53.9 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
12|1500 A              | 1.04      ||microJy             |2.00E+15|  1.04E-06||Jy|2010ApJ...723..241S|no uncertainty reported|      1500 A         | Broad-band measurement|12 36 45.71 +62 07 54.3 (J2000)| Flux in fixed aperture|                                        |Transformed from previously published data;Extinction-corrected for Milky Way
13|u (SDSS PSF) AB     | 22.895    |+/-0.448|asinh mag           |8.36E+14|  2.51E-06|+/-1.12E-06|Jy|2007SDSS6.C...0000:|based on count statistics only|3585       A         | Broad-band measurement|189.1905450554 62.1317861452 (J2000)| Modelled datum|SDSS flags: CANONICAL_CENTER - used canonical, not local, center; NOPETRO - no Petrosian radius could be determined; MANYR90 - more than one 90% radius; BAD_RADIAL - some low S/N radial points; PETROFAINT - Petrosian radius measured at very low surface brightness; ELLIPFAINT - no isophotal fits performed; AMOMENT_FAINT - too faint for adaptive moments;|From new raw data
14|U (KPNO) AB         | 23.6      || mag                |8.22E+14|  1.32E-06||Jy|2004AJ....127.3137C|no uncertainty reported| 3647.65   A         | Broad-band measurement|189.190475 +62.13182 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
15|B F435W (HST/ACS) AB      | 23.487    ||mag                 |6.98E+14|  1.46E-06||Jy|2007ApJ...660...81M|no uncertainty reported|    4297   A         | Broad-band measurement|12 36 45.783 +62 07 54.27 (J2000)| Flux integrated from map|                                        |From reprocessed raw data; Corrected for contaminatingsources
16|B (Subaru) AB       | 23.39     ||mag                 |6.77E+14|  1.60E-06||Jy|2006ApJ...653.1027W|no uncertainty reported| 4427.60   A         | Broad-band measurement|189.190763 62.131742 (J2000)| Flux in fixed aperture|3" diameter aperture                    |Averaged from previously published data
17|B (Subaru) AB       | 23.4      || mag                |6.77E+14|  1.59E-06||Jy|2004AJ....127.3137C|no uncertainty reported| 4427.60   A         | Broad-band measurement|189.190475 +62.13182 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
18|g (SDSS PSF) AB     | 23.542    |+/-0.295|asinh mag           |6.17E+14|  1.31E-06|+/-3.99E-07|Jy|2007SDSS6.C...0000:|based on count statistics only|4858       A         | Broad-band measurement|189.1905450554 62.1317861452 (J2000)| Modelled datum|SDSS flags: CANONICAL_CENTER - used canonical, not local, center; NOPETRO - no Petrosian radius could be determined; BAD_RADIAL - some low S/N radial points; PETROFAINT - Petrosian radius measured at very low surface brightness; ELLIPFAINT - no isophotal fits performed; AMOMENT_FAINT - too faint for adaptive moments;|From new raw data
19|V (Subaru) AB       | 23.4      || mag                |5.48E+14|  1.59E-06||Jy|2004AJ....127.3137C|no uncertainty reported| 5471.22   A         | Broad-band measurement|189.190475 +62.13182 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
20|V (HST/ACS) AB      | 23.222    ||mag                 |5.08E+14|  1.87E-06||Jy|2007ApJ...660...81M|no uncertainty reported|    5907   A         | Broad-band measurement|12 36 45.783 +62 07 54.27 (J2000)| Flux integrated from map|                                        |From reprocessed raw data; Corrected for contaminatingsources
21|r (SDSS PSF) AB     | 22.618    |+/-0.192|asinh mag           |4.77E+14|  3.20E-06|+/-5.86E-07|Jy|2007SDSS6.C...0000:|based on count statistics only|6290       A         | Broad-band measurement|189.1905450554 62.1317861452 (J2000)| Modelled datum|SDSS flags: NOPETRO - no Petrosian radius could be determined; BAD_RADIAL - some low S/N radial points; PETROFAINT - Petrosian radius measured at very low surface brightness; ELLIPFAINT - no isophotal fits performed; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding; CANONICAL_BAND - this band was primary (usually r);|From new raw data
22|R (Keck II) AB      | 23.00     || mag                |4.62E+14|  2.29E-06||Jy|2004AJ....127.3121W|no uncertainty reported|   648.7   A         | Broad-band measurement|12 36 45.783 +62 07 54.27 (J2000)| Total flux|                                        |From new raw data
23|R (Subaru) AB       | 22.89     ||mag                 |4.59E+14|  2.54E-06||Jy|2006ApJ...653.1027W|no uncertainty reported| 6534.16   A         | Broad-band measurement|189.190763 62.131742 (J2000)| Flux in fixed aperture|3" diameter aperture                    |Averaged from previously published data
24|R (Subaru) AB       | 22.9      || mag                |4.59E+14|  2.51E-06||Jy|2004AJ....127.3137C|no uncertainty reported| 6534.16   A         | Broad-band measurement|189.190475 +62.13182 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
25|i (SDSS PSF) AB     | 22.211    |+/-0.238|asinh mag           |3.89E+14|  4.65E-06|+/-1.06E-06|Jy|2007SDSS6.C...0000:|based on count statistics only|7706       A         | Broad-band measurement|189.1905450554 62.1317861452 (J2000)| Modelled datum|SDSS flags: CANONICAL_CENTER - used canonical, not local, center; BAD_RADIAL - some low S/N radial points; INTERP - object contains interpolated-over pixels; ELLIPFAINT - no isophotal fits performed;|From new raw data
26|i F775W (HST/ACS) AB      | 22.837    ||mag                 |3.86E+14|  2.66E-06||Jy|2007ApJ...660...81M|no uncertainty reported|    7764   A         | Broad-band measurement|12 36 45.783 +62 07 54.27 (J2000)| Flux integrated from map|                                        |From reprocessed raw data; Corrected for contaminatingsources
27|I (Subaru) AB       | 22.6      || mag                |3.76E+14|  3.31E-06||Jy|2004AJ....127.3137C|no uncertainty reported| 7975.89   A         | Broad-band measurement|189.190475 +62.13182 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
28|I (Subaru) AB       | 22.56     ||mag                 |3.76E+14|  3.44E-06||Jy|2006ApJ...653.1027W|no uncertainty reported| 7975.89   A         | Broad-band measurement|189.190763 62.131742 (J2000)| Flux in fixed aperture|3" diameter aperture                    |Averaged from previously published data
29|z' (Subaru) AB      | 22.2      || mag                |3.31E+14|  4.79E-06||Jy|2004AJ....127.3137C|no uncertainty reported| 9069.21   A         | Broad-band measurement|189.190475 +62.13182 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
30|z (SDSS PSF) AB     | 21.224    |+/-0.402|asinh mag           |3.25E+14|  1.09E-05|+/-4.50E-06|Jy|2007SDSS6.C...0000:|based on count statistics only|9222       A         | Broad-band measurement|189.1905450554 62.1317861452 (J2000)| Modelled datum|SDSS flags: CANONICAL_CENTER - used canonical, not local, center; BAD_RADIAL - some low S/N radial points; ELLIPFAINT - no isophotal fits performed; AMOMENT_FAINT - too faint for adaptive moments;|From new raw data
31|z F850LP (HST/ACS) AB      | 22.288    ||mag                 |3.17E+14|  4.41E-06||Jy|2007ApJ...660...81M|no uncertainty reported|    9445   A         | Broad-band measurement|12 36 45.783 +62 07 54.27 (J2000)| Flux integrated from map|                                        |From reprocessed raw data; Corrected for contaminatingsources
32|HK' (QUIRC) AB      | 20.90     |+/-0.15 |mag                 |1.58E+14|  1.59E-05|+/-2.19E-06|Jy|2006ApJ...653.1027W|uncertainty|18947.38   A         | Broad-band measurement|189.190763 62.131742 (J2000)| Flux in fixed aperture|3" diameter aperture                    |Averaged from previously published data
33|HK' (UH) AB         | 20.9      || mag                |1.58E+14|  1.59E-05||Jy|2004AJ....127.3137C|no uncertainty reported|18947.38   A         | Broad-band measurement|189.190475 +62.13182 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
34|3.6 microns (IRAC)  | 38.20     |+/-1.91 |microJy             |8.44E+13|  3.82E-05|+/-1.91E-06|Jy|2011AJ....141....1T|rms uncertainty|     3.550 microns   | Broad-band measurement|189.190948 62.131733 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
35|4.5 microns (IRAC)  | 44.00     |+/-2.20 |microJy             |6.67E+13|  4.40E-05|+/-2.20E-06|Jy|2011AJ....141....1T|rms uncertainty|     4.493 microns   | Broad-band measurement|189.190948 62.131733 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
36|5.8 microns (IRAC)  | 34.80     |+/-1.80 |microJy             |5.23E+13|  3.48E-05|+/-1.80E-06|Jy|2011AJ....141....1T|rms uncertainty|     5.731 microns   | Broad-band measurement|189.190948 62.131733 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
37|8.0 microns (IRAC)  | 44.80     |+/-2.31 |microJy             |3.81E+13|  4.48E-05|+/-2.31E-06|Jy|2011AJ....141....1T|rms uncertainty|     7.872 microns   | Broad-band measurement|189.190948 62.131733 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
38|16 microns (IRS)    | 323.4     |+/-15.2 |microJy             |1.90E+13|  3.23E-04|+/-1.52E-05|Jy|2011AJ....141....1T|rms uncertainty|      15.8 microns   | Broad-band measurement|189.190948 62.131733 (J2000)| From fitting to map|                                        |From new raw data
39|24 microns (MIPS)   | 374.0     |+/-7.9  |microJy             |1.27E+13|  3.74E-04|+/-7.90E-06|Jy|2011AJ....141....1T|rms uncertainty|     23.68 microns   | Broad-band measurement|189.190948 62.131733 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
1|24 microns (MIPS)   | 0.172     |+/-0.034|mJy             |1.27E+13|172.E-06|+/-34.0E-06|Jy|2009ApJ...694.1517D|3sigma uncertainty|     23.68 microns   | Broad-band measurement|12 37 11.89 +62 22 11.8 (J2000)| Flux integrated from map|                                        |From new raw data
40|24 microns (MIPS)   | 369       |+/-7    |microJy             |1.27E+13|  3.69E-04|+/-7.00E-06|Jy|2011ApJ...726...93R|uncertainty|     23.68 microns   | Broad-band measurement|12 36 45.89 +62 07 54.1 (J2000)| Not reported in paper|                                        |Averaged from previously published data
2|24 microns (MIPS)   | 0.366     |+/-0.006|mJy             |1.27E+13|0.366E-03|+/-0.006E-03|Jy|2009ApJ...694.1517D|3sigma uncertainty|     23.68 microns   | Broad-band measurement|12 37 11.89 +62 22 11.8 (J2000)| Flux integrated from map|                                        |From new raw data
41|24 microns (MIPS)   | 371.4     |+/-5.0  |microJy             |1.27E+13|  3.71E-04|+/-5.00E-06|Jy|2011A&A...528A..35M|uncertainty|     23.68 microns   | Broad-band measurement|12 36 45.83 +62 07 54.17 (J2000)| Flux integrated from map|                                        |From new raw data
42|70 microns (MIPS)   | 4.8       |+/-0.4  | milliJy            |4.20E+12|  4.80E-03|+/-4.00E-04|Jy|2009MNRAS.399..121C|uncertainty|     71.42 microns   | Broad-band measurement|123645.89 +620754.1 (J2000)| Flux integrated from map|                                        |From reprocessed raw data
43|70 microns (MIPS)   | 6.1       |+/-0.4  |milliJy             |4.20E+12|  6.10E-03|+/-4.00E-04|Jy|2011A&A...528A..35M|uncertainty|     71.42 microns   | Broad-band measurement|12 36 45.83 +62 07 54.17 (J2000)| Flux integrated from map|                                        |From new raw data
4|70 microns (MIPS)   | 5.6       |+/-0.7  |mJy             |4.20E+12|5.6E-03 |+/-0.7E-03|Jy|2009ApJ...699.1610H|3 sigma|     71.42 microns   | Broad-band measurement|221804.42 +002154.4 (J2000)| Flux in fixed aperture|                                        |From new raw data
44|850 microns (SCUBA) ||<6.3       | milliJy            |3.53E+11||6.30E-03|Jy|2009MNRAS.399..121C|2 sigma|       850 microns   | Broad-band measurement|123645.89 +620754.1 (J2000)| Flux integrated from map|                                        |From new raw data
5|850 microns (SCUBA) |           |<16.2   |mJy             |3.53E+11|        |16.2E-03|Jy|2005MNRAS.358..149P|3rms uncertainty|     850   microns   | Broad-band measurement|12 37 11.7 +62 22 12 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
6|1200 microns (MAMBO)|           |<2.4    |mJy             |2.50E+11|        |2.4E-03|Jy|2004MNRAS.354..779G|3rms uncertainty|      1200 microns   | Broad-band measurement|16 36 55.9 +40 59 12 (J2000)| Flux integrated from map|S/N = 3.66                              |From new raw data
45|1.4 GHz (MERLIN)    | 83.4      |+/-9.8  | microJy            |1.40E+09|  8.34E-05|+/-9.80E-06|Jy|2009MNRAS.399..121C|uncertainty|       1.4 GHz       | Broad-band measurement|123645.89 +620754.1 (J2000)| Flux integrated from map|                                        |From new raw data
46|1.4 GHz (VLA)       | 73.2      |+/-5.6  |microJy             |1.40E+09|  7.32E-05|+/-5.60E-06|Jy|2010ApJS..188..178M|uncertainty|       1.4 GHz       | Broad-band measurement|12 36 45.82 +62 07 54.3 (J2000)| Total flux; Beam filling or dilution corrected|Major=2.0"; Minor=0.0"; PA=80 deg       |From new raw data
47|1.4 GHz (VLA)       | 49        ||microJy             |1.40E+09|  4.90E-05||Jy|2005MNRAS.358.1159M|no uncertainty reported|     1.4   GHz       | Broad-band measurement|12 36 45.862 +62 07 54.19 (J2000)| Flux integrated from map|                                        |From new raw data
48|1.4 GHz             | 48.9      |+/-8.4  |microJy             |1.40E+09|  4.89E-05|+/-8.40E-06|Jy|2000ApJ...533..611R|1 sigma|1.4        GHz       | Broad-band measurement; broad-band flux derived by integration over spectrum; synthetic band|123645.875 +620754.25 (J2000)| Flux integrated from map; Pointing and beam filling|                                        |From new raw data; Corrected for contaminating sources
49|1.4 GHz (VLA)       | 66        |+/-12   | microJy            |1.40E+09|  6.60E-05|+/-1.20E-05|Jy|2006MNRAS.371..963B|1 sigma|       1.4 GHz       | Broad-band measurement|12 36 45.827 +62 07 54.26 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
