
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-07-10T02:51:09PDT



Photometric Data for SDSS J091127.61+055054.0

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|2-10 keV (XMM)      | 1.8E-13   || erg/cm^2^/s        |1.45E+18|  1.24E-08||Jy|2009ApJS..183...17Y|no uncertainty reported|      6.00 keV       | Broad-band measurement|091127.61 +055054.0 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
2|2-10 keV (XMM)      | -12.80    ||log(erg/s/cm^2^)    |1.45E+18|  1.09E-08||Jy|2010A&A...515A...2S|no uncertainty reported|      6.00 keV       | Broad-band measurement|| Modelled datum|                                        |From reprocessed raw data; NED frequency assigned tomid-point of band in keV
3|2-10 keV (XMM)      | -12.8     ||log(erg/s/cm^2^)    |1.45E+18|  1.09E-08||Jy|2008A&A...491..425G|no uncertainty reported|      6.00 keV       | Broad-band measurement|| Modelled datum|                                        |From reprocessed raw data; Extinction-corrected for MilkyWay; NED frequency assigned to mid-point of band in keV
4|0.3-10 keV (XMM)    | 0.2E-12   ||erg cm^-2^ s^-1^    |1.25E+18|  1.60E-08||Jy|2005MNRAS.364..195P|no uncertainty reported|    5.15   keV       | Broad-band measurement|09 11 27.5 +05 50 52.0 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
5|0.3-10 keV (XMM)    | -12.620   || log(erg/cm^2^/s)   |1.25E+18|  1.92E-08||Jy|2009ApJ...690.1006F|no uncertainty reported|      5.15 keV       | Broad-band measurement|091127.61 +055054.1 (J2000)| Flux integrated from map|                                        |From reprocessed raw data; NED frequency assigned tomid-point of band in keV
6|0.5-8 keV (Chandra) | 1.9E-14   |+/-0.8E-14|ergs/cm^2^/s        |1.03E+18|  1.84E-09|+/-7.77E-10|Jy|2007ApJ...661...19P|uncertainty|    4.25   keV       | Broad-band measurement|| From fitting to map|Unabsorbed flux                         |From reprocessed raw data; NED frequency assigned tomid-point of band in keV
7|0.5-8 keV (Chandra) | 1.8E-14   |+/-0.5E-14|ergs/cm^2^/s        |1.03E+18|  1.75E-09|+/-4.85E-10|Jy|2007ApJ...661...19P|uncertainty|    4.25   keV       | Broad-band measurement|| From fitting to map|Unabsorbed flux                         |From reprocessed raw data; NED frequency assigned tomid-point of band in keV
8|0.5-8 keV (Chandra) | 1.24E-13  |+/-0.99E-13|erg/cm^2^/s         |1.03E+18|  1.20E-08|+/-9.61E-09|Jy|2012ApJ...744..111P|uncertainty|      4.25 keV       | Broad-band measurement|| Total flux|                                        |From reprocessed raw data; Extinction-corrected for MilkyWay; NED frequency assigned to mid-point of band in keV
9|0.4-8 keV (Chandra) | 1.1E-13   ||ergs/cm^2^/s        |1.02E+18|  1.08E-08||Jy|2004ApJ...605...45D|no uncertainty reported|    4.20   keV       | Broad-band measurement|| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
10|0.5-2 keV (XMM)     | 4.0E-14   || erg/cm^2^/s        |3.02E+17|  1.32E-08||Jy|2009ApJS..183...17Y|no uncertainty reported|      1.25 keV       | Broad-band measurement|091127.61 +055054.0 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
11|0.5-2 keV (XMM)     | -13.29    ||log(erg/s/cm^2^)    |3.02E+17|  1.70E-08||Jy|2010A&A...515A...2S|no uncertainty reported|      1.25 keV       | Broad-band measurement|| Modelled datum|                                        |From reprocessed raw data; NED frequency assigned tomid-point of band in keV
12|0.5-2 keV (XMM)     | -13.3     ||log(erg/s/cm^2^)    |3.02E+17|  1.66E-08||Jy|2008A&A...491..425G|no uncertainty reported|      1.25 keV       | Broad-band measurement|| Modelled datum|                                        |From reprocessed raw data; Extinction-corrected for MilkyWay; NED frequency assigned to mid-point of band in keV
13|FUV (GALEX)         | 28.248E-17|| erg/s/cm^2^/A      |1.98E+15|  2.17E-05||Jy|2009ApJ...690.1181S|no uncertainty reported|      1516 A         | Broad-band measurement|137.865070 +05.848365 (J2000)| Not reported in paper|                                        |Averaged from previously published data
14|FUV (GALEX)         | 18.94E-17 ||erg/s/cm^2^/A       |1.95E+15|  1.50E-05||Jy|2009ApJS..185...20S|no uncertainty reported|      1539 A         | Broad-band measurement|137.865067 +05.84835 (J2000)| Flux in fixed aperture|                                        |Transformed from previously published data
15|1700 A (SDSS)       | -15.128   ||log(erg/cm^2^/s/A)  |1.76E+15|  7.19E-05||Jy|2011MNRAS.410..860A|no uncertainty reported|      1700 A         | Broad-band measurement|137.865067 +05.848365 (J2000)| Flux integrated from map|                                        |From reprocessed raw data
16|NUV (GALEX)         | 28.355E-17|| erg/s/cm^2^/A      |1.32E+15|  4.87E-05||Jy|2009ApJ...690.1181S|no uncertainty reported|      2267 A         | Broad-band measurement|137.865070 +05.848365 (J2000)| Not reported in paper|                                        |Averaged from previously published data
17|NUV (GALEX)         | 22.87E-17 ||erg/s/cm^2^/A       |1.29E+15|  4.10E-05||Jy|2009ApJS..185...20S|no uncertainty reported|      2316 A         | Broad-band measurement|137.865067 +05.84835 (J2000)| Flux in fixed aperture|                                        |Transformed from previously published data
18|u (SDSS PSF) AB     | 18.890    |+/-0.027|asinh mag           |8.36E+14|  1.05E-04|+/-2.60E-06|Jy|2007SDSS6.C...0000:|based on count statistics only|3585       A         | Broad-band measurement|137.8650599181 5.8483668713 (J2000)| Modelled datum|SDSS flags: CHILD - object is part of a blended parent object; BAD_RADIAL - some low S/N radial points; INTERP - object contains interpolated-over pixels; BINNED1 - detected at >=5 sigma in original imaging frame;|From new raw data
19|u (SDSS Model) AB   | 18.799    |+/-0.021|asinh mag           |8.36E+14|  1.14E-04|+/-2.16E-06|Jy|2004SDSS3.C...0000:|based on count statistics only|3585       A         | Broad-band measurement|137.865051 5.848367 (J2000)| Modelled datum|SDSS flags: CHILD - object is part of a blended parent object; BAD_RADIAL - some low S/N radial points; INTERP - object contains interpolated-over pixels; BINNED1 - detected at >=5 sigma in original imaging frame;|From new raw data
20|u (SDSS PSF) AB     | 18.890    |+/-0.027|asinh mag           |8.36E+14|  1.05E-04|+/-2.58E-06|Jy|2004SDSS3.C...0000:|based on count statistics only|3585       A         | Broad-band measurement|137.865051 5.848367 (J2000)| Modelled datum|SDSS flags: CHILD - object is part of a blended parent object; BAD_RADIAL - some low S/N radial points; INTERP - object contains interpolated-over pixels; BINNED1 - detected at >=5 sigma in original imaging frame;|From new raw data
21|u (SDSS Petrosian)AB| 18.850    |+/-0.030|asinh mag           |8.36E+14|  1.09E-04|+/-3.00E-06|Jy|2004SDSS3.C...0000:|based on count statistics only|3585       A         | Broad-band measurement|137.865051 5.848367 (J2000)| Modelled datum|From new raw data
22|u (SDSS CModel) AB  | 18.790    ||asinh mag           |8.36E+14|  1.11E-04||Jy|2004SDSS3.C...0000:|no uncertainty reported|3585       A         | Broad-band measurement|137.865051 5.848367 (J2000)| Modelled datum|SDSS flags: CHILD - object is part of a blended parent object; BAD_RADIAL - some low S/N radial points; INTERP - object contains interpolated-over pixels; BINNED1 - detected at >=5 sigma in original imaging frame;|From new raw data
23|g (SDSS PSF) AB     | 18.023    |+/-0.026|asinh mag           |6.17E+14|  2.24E-04|+/-5.37E-06|Jy|2007SDSS6.C...0000:|based on count statistics only|4858       A         | Broad-band measurement|137.8650599181 5.8483668713 (J2000)| Modelled datum|SDSS flags: CHILD - object is part of a blended parent object; BAD_RADIAL - some low S/N radial points; BINNED1 - detected at >=5 sigma in original imaging frame;|From new raw data
24|g (SDSS CModel) AB  | 17.937    ||asinh mag           |6.17E+14|  2.43E-04||Jy|2004SDSS3.C...0000:|no uncertainty reported|4858       A         | Broad-band measurement|137.865051 5.848367 (J2000)| Modelled datum|SDSS flags: CHILD - object is part of a blended parent object; BAD_RADIAL - some low S/N radial points; BINNED1 - detected at >=5 sigma in original imaging frame;|From new raw data
25|g (SDSS Model) AB   | 17.940    |+/-0.006|asinh mag           |6.17E+14|  2.42E-04|+/-1.30E-06|Jy|2004SDSS3.C...0000:|based on count statistics only|4858       A         | Broad-band measurement|137.865051 5.848367 (J2000)| Modelled datum|SDSS flags: CHILD - object is part of a blended parent object; BAD_RADIAL - some low S/N radial points; BINNED1 - detected at >=5 sigma in original imaging frame;|From new raw data
26|g (SDSS Petrosian)AB| 17.991    |+/-0.012|asinh mag           |6.17E+14|  2.31E-04|+/-2.58E-06|Jy|2004SDSS3.C...0000:|based on count statistics only|4858       A         | Broad-band measurement|137.865051 5.848367 (J2000)| Modelled datum|From new raw data
27|g (SDSS PSF) AB     | 18.023    |+/-0.026|asinh mag           |6.17E+14|  2.24E-04|+/-5.33E-06|Jy|2004SDSS3.C...0000:|based on count statistics only|4858       A         | Broad-band measurement|137.865051 5.848367 (J2000)| Modelled datum|SDSS flags: CHILD - object is part of a blended parent object; BAD_RADIAL - some low S/N radial points; BINNED1 - detected at >=5 sigma in original imaging frame;|From new raw data
28|F555W (HST/WFPC2)         | 22.97     |+/-0.22 | mag                |5.54E+14|  2.42E-06|+/-4.90E-07|Jy|2008A&A...478...95Y|uncertainty|      5407 A         | Broad-band measurement|| Modelled datum|                                        |Averaged from previously published data
29|r (SDSS Petrosian)AB| 17.824    |+/-0.014|asinh mag           |4.77E+14|  2.69E-04|+/-3.49E-06|Jy|2004SDSS3.C...0000:|based on count statistics only|6290       A         | Broad-band measurement|137.865051 5.848367 (J2000)| Modelled datum|From new raw data
30|r (SDSS PSF) AB     | 17.884    |+/-0.018|asinh mag           |4.77E+14|  2.55E-04|+/-4.20E-06|Jy|2004SDSS3.C...0000:|based on count statistics only|6290       A         | Broad-band measurement|137.865051 5.848367 (J2000)| Modelled datum|SDSS flags: CHILD - object is part of a blended parent object; BAD_RADIAL - some low S/N radial points; BINNED1 - detected at >=5 sigma in original imaging frame; CANONICAL_BAND - this band was primary (usually r);|From new raw data
31|r (SDSS PSF) AB     | 17.884    |+/-0.018|asinh mag           |4.77E+14|  2.55E-04|+/-4.23E-06|Jy|2007SDSS6.C...0000:|based on count statistics only|6290       A         | Broad-band measurement|137.8650599181 5.8483668713 (J2000)| Modelled datum|SDSS flags: CHILD - object is part of a blended parent object; BAD_RADIAL - some low S/N radial points; BINNED1 - detected at >=5 sigma in original imaging frame; CANONICAL_BAND - this band was primary (usually r);|From new raw data
32|r (SDSS CModel) AB  | 17.778    ||asinh mag           |4.77E+14|  2.81E-04||Jy|2004SDSS3.C...0000:|no uncertainty reported|6290       A         | Broad-band measurement|137.865051 5.848367 (J2000)| Modelled datum|SDSS flags: CHILD - object is part of a blended parent object; BAD_RADIAL - some low S/N radial points; BINNED1 - detected at >=5 sigma in original imaging frame; CANONICAL_BAND - this band was primary (usually r);|From new raw data
33|r (SDSS Model) AB   | 17.778    |+/-0.006|asinh mag           |4.77E+14|  2.81E-04|+/-1.57E-06|Jy|2004SDSS3.C...0000:|based on count statistics only|6290       A         | Broad-band measurement|137.865051 5.848367 (J2000)| Modelled datum|SDSS Effective Radius =   0.13" x   0.06".;SDSS flags: CHILD - object is part of a blended parent object; BAD_RADIAL - some low S/N radial points; BINNED1 - detected at >=5 sigma in original imaging frame; CANONICAL_BAND - this band was primary (usually r);|From new raw data
34|i (SDSS Model) AB   | 17.765    |+/-0.008|asinh mag           |3.89E+14|  2.84E-04|+/-1.97E-06|Jy|2004SDSS3.C...0000:|based on count statistics only|7706       A         | Broad-band measurement|137.865051 5.848367 (J2000)| Modelled datum|SDSS flags: CHILD - object is part of a blended parent object; BAD_RADIAL - some low S/N radial points; BINNED1 - detected at >=5 sigma in original imaging frame; BRIGHTEST_GALAXY_CHILD - brightest child among one parent's children;|From new raw data
35|i (SDSS PSF) AB     | 17.911    |+/-0.020|asinh mag           |3.89E+14|  2.49E-04|+/-4.65E-06|Jy|2004SDSS3.C...0000:|based on count statistics only|7706       A         | Broad-band measurement|137.865051 5.848367 (J2000)| Modelled datum|SDSS flags: CHILD - object is part of a blended parent object; BAD_RADIAL - some low S/N radial points; BINNED1 - detected at >=5 sigma in original imaging frame; BRIGHTEST_GALAXY_CHILD - brightest child among one parent's children;|From new raw data
36|i (SDSS Petrosian)AB| 17.771    |+/-0.015|asinh mag           |3.89E+14|  5.75E-04|+/-8.16E-06|Jy|2004SDSS3.C...0000:|based on count statistics only|7706       A         | Broad-band measurement|137.865051 5.848367 (J2000)| Modelled datum|From new raw data
37|i (SDSS CModel) AB  | 17.751    ||asinh mag           |3.89E+14|  2.88E-04||Jy|2004SDSS3.C...0000:|no uncertainty reported|7706       A         | Broad-band measurement|137.865051 5.848367 (J2000)| Modelled datum|SDSS flags: CHILD - object is part of a blended parent object; BAD_RADIAL - some low S/N radial points; BINNED1 - detected at >=5 sigma in original imaging frame; BRIGHTEST_GALAXY_CHILD - brightest child among one parent's children;|From new raw data
38|i (SDSS PSF) AB     | 17.911    |+/-0.020|asinh mag           |3.89E+14|  2.49E-04|+/-4.58E-06|Jy|2007SDSS6.C...0000:|based on count statistics only|7706       A         | Broad-band measurement|137.8650599181 5.8483668713 (J2000)| Modelled datum|SDSS flags: CHILD - object is part of a blended parent object; BAD_RADIAL - some low S/N radial points; BINNED1 - detected at >=5 sigma in original imaging frame; BRIGHTEST_GALAXY_CHILD - brightest child among one parent's children;|From new raw data
39|F814W (HST/WFPC2)         | 20.47     |+/-0.09 | mag                |3.78E+14|  1.62E-05|+/-1.34E-06|Jy|2008A&A...478...95Y|uncertainty|      7940 A         | Broad-band measurement|| Modelled datum|                                        |Averaged from previously published data
40|I (HST)             | 17.39     ||mag                 |3.68E+14|  2.67E-04||Jy|2011ApJ...738...96M|no uncertainty reported|     0.814 microns   | Broad-band measurement|| Not reported in paper|                                        |From reprocessed raw data
41|z (SDSS Petrosian)AB| 17.852    |+/-0.038|asinh mag           |3.25E+14|  2.58E-04|+/-8.97E-06|Jy|2004SDSS3.C...0000:|based on count statistics only|9222       A         | Broad-band measurement|137.865051 5.848367 (J2000)| Modelled datum|From new raw data
42|z (SDSS PSF) AB     | 17.895    |+/-0.027|asinh mag           |3.25E+14|  2.48E-04|+/-6.27E-06|Jy|2004SDSS3.C...0000:|based on count statistics only|9222       A         | Broad-band measurement|137.865051 5.848367 (J2000)| Modelled datum|SDSS flags: CHILD - object is part of a blended parent object; BAD_RADIAL - some low S/N radial points; BINNED1 - detected at >=5 sigma in original imaging frame;|From new raw data
43|z (SDSS CModel) AB  | 17.756    ||asinh mag           |3.25E+14|  2.87E-04||Jy|2004SDSS3.C...0000:|no uncertainty reported|9222       A         | Broad-band measurement|137.865051 5.848367 (J2000)| Modelled datum|SDSS flags: CHILD - object is part of a blended parent object; BAD_RADIAL - some low S/N radial points; BINNED1 - detected at >=5 sigma in original imaging frame;|From new raw data
44|z (SDSS Model) AB   | 17.781    |+/-0.020|asinh mag           |3.25E+14|  2.75E-04|+/-4.95E-06|Jy|2004SDSS3.C...0000:|based on count statistics only|9222       A         | Broad-band measurement|137.865051 5.848367 (J2000)| Modelled datum|SDSS flags: CHILD - object is part of a blended parent object; BAD_RADIAL - some low S/N radial points; BINNED1 - detected at >=5 sigma in original imaging frame;|From new raw data
45|z (SDSS PSF) AB     | 17.895    |+/-0.027|asinh mag           |3.25E+14|  2.48E-04|+/-6.16E-06|Jy|2007SDSS6.C...0000:|based on count statistics only|9222       A         | Broad-band measurement|137.8650599181 5.8483668713 (J2000)| Modelled datum|SDSS flags: CHILD - object is part of a blended parent object; BAD_RADIAL - some low S/N radial points; BINNED1 - detected at >=5 sigma in original imaging frame;|From new raw data
46|F160W (HST/NICMOS)         | 17.93     |+/-0.08 | mag                |1.87E+14|  7.02E-05|+/-5.17E-06|Jy|2008A&A...478...95Y|uncertainty|     1.603 microns   | Broad-band measurement|| Modelled datum|                                        |Averaged from previously published data
47|350 microns (CSO/SHARC-II)   | 150       |+/-21   |milliJy             |8.57E+11|  1.50E-01|+/-2.10E-02|Jy|2009ApJ...707..988W|rms noise|       350 microns   | Broad-band measurement|09 11 27.40 +05 50 52.0 (J2000)| Flux integrated from map|S/N=7.1 sigma                           |From new raw data
3|450 microns (SCUBA) | 65.0 |+/-19.0      | milliJy            |6.66E+11| 65.E-3|19.E-3|Jy|2008MNRAS.384.1611K| uncertainty reported|       450 microns   | Broad-band measurement|163555.5 +661300 (J2000)| Flux integrated from map|                                        |From new raw data
5|850 microns (SCUBA) | 26.7      |+/-1.4  | milliJy            |3.53E+11|  26.7E-03|+/-1.40E-03|Jy|2008MNRAS.384.1611K|rms uncertainty|       850 microns   | Broad-band measurement|163555.5 +661300 (J2000)| Flux integrated from map|S/N = 15.8                              |From new raw data
48|CO(3-2) (OVRO)      | 2.9       |+/-1.1  | Jy km/s            |3.46E+11|  8.81E+05|+/-3.34E+05|Jy-Hz|2004ApJ...609...61H|uncertainty|   2.796             | Line measurement; flux integrated over line; lines measured in emission|09 11 27.50 +05 50 52.0 (J2000)| Flux integrated from map|                                        |From new raw data
27|1.3 mm (PdBI)       | 10.2       |+/-1.8  |milliJy             |2.31E+11|  10.2E-03|+/-1.8E-03|Jy|2006ApJ...640..228T|uncertainty|     1.3   mm        | Broad-band measurement| | Flux integrated from map|                                        |From new raw data
49|CO(1-0) (EVLA)      | 0.205     |+/-0.029|Jy km/s             |1.15E+11|  2.08E+04|+/-2.94E+03|Jy-Hz|2011ApJ...739L..32R|uncertainty|   115.271 GHz       | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|                                        |From new raw data
9|100.8 GHz (IRAM/PdBI) | 1.7       |+/-0.3  | milliJy            |1.008E+11|  1.7E-03|+/-0.3E-03|Jy|2007A&A...470...53A|uncertainty|       110 GHz       | Broad-band measurement|| From fitting to map|                                        |From new raw data
