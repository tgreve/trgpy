
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2017-01-17T08:25:23PST



Photometric Data for Cosmic Eyelash

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|F336W (HST/ACS)         ||<0.1       |microJy             |8.97E+14||1.00E-07|Jy|2010Natur.464..733S|no uncertainty reported|      3344 A         | Broad-band measurement|21 35 11.6 -01 02 52.0 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
2|F606W (HST/ACS)         | 0.9       |+/-0.2  |microJy             |5.08E+14|  9.00E-07|+/-2.00E-07|Jy|2010Natur.464..733S|uncertainty|      5907 A         | Broad-band measurement|21 35 11.6 -01 02 52.0 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
3|F814W (HST/ACS)         | 1.4       |+/-0.4  |microJy             |3.74E+14|  1.40E-06|+/-4.00E-07|Jy|2010Natur.464..733S|uncertainty|      8012 A         | Broad-band measurement|21 35 11.6 -01 02 52.0 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
4|K (UKIRT)           | 36        |+/-4    |microJy             |1.37E+14|  3.60E-05|+/-4.00E-06|Jy|2010Natur.464..733S|uncertainty|     2.195 microns   | Broad-band measurement|21 35 11.6 -01 02 52.0 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
5|3.6 microns (IRAC)  | 1.5495E+02|+/-8.2675E-01|microJy             |8.44E+13|  1.55E-04|+/-8.27E-07|Jy|2013SSTSLC4.2....0C|uncertainty|3.55       microns   | Broad-band measurement|| Flux in fixed aperture|5.8" aperture                           |From new raw data
6|3.6 microns (IRAC)  | 8.2719E+01|+/-5.8968E-01|microJy             |8.44E+13|  8.27E-05|+/-5.90E-07|Jy|2013SSTSLC4.2....0C|uncertainty|3.55       microns   | Broad-band measurement|| Flux in fixed aperture|3.8" aperture                           |From new raw data
7|3.6 microns (IRAC)  | 0.13      |+/-0.02 |milliJy             |8.44E+13|  1.30E-04|+/-2.00E-05|Jy|2010Natur.464..733S|uncertainty|     3.550 microns   | Broad-band measurement|21 35 11.6 -01 02 52.0 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
8|4.5 microns (IRAC)  | 1.4681E+02|+/-1.0325E+00|microJy             |6.67E+13|  1.47E-04|+/-1.03E-06|Jy|2013SSTSLC4.2....0C|uncertainty|4.493      microns   | Broad-band measurement|| Flux in fixed aperture|3.8" aperture                           |From new raw data
9|4.5 microns (IRAC)  | 2.3641E+02|+/-1.3766E+00|microJy             |6.67E+13|  2.36E-04|+/-1.38E-06|Jy|2013SSTSLC4.2....0C|uncertainty|4.493      microns   | Broad-band measurement|| Flux in fixed aperture|5.8" aperture                           |From new raw data
10|4.5 microns (IRAC)  | 0.21      |+/-0.02 |milliJy             |6.67E+13|  2.10E-04|+/-2.00E-05|Jy|2010Natur.464..733S|uncertainty|     4.493 microns   | Broad-band measurement|21 35 11.6 -01 02 52.0 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
11|5.8 microns (IRAC)  | 3.5479E+02|+/-3.9105E+00|microJy             |5.23E+13|  3.55E-04|+/-3.91E-06|Jy|2013SSTSLC4.2....0C|uncertainty|5.731      microns   | Broad-band measurement|| Flux in fixed aperture|5.8" aperture                           |From new raw data
12|5.8 microns (IRAC)  | 2.7517E+02|+/-3.3566E+00|microJy             |5.23E+13|  2.75E-04|+/-3.36E-06|Jy|2013SSTSLC4.2....0C|uncertainty|5.731      microns   | Broad-band measurement|| Flux in fixed aperture|3.8" aperture                           |From new raw data
13|5.8 microns (IRAC)  | 0.32      |+/-0.05 |milliJy             |5.23E+13|  3.20E-04|+/-5.00E-05|Jy|2010Natur.464..733S|uncertainty|     5.731 microns   | Broad-band measurement|21 35 11.6 -01 02 52.0 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
14|8.0 microns (IRAC)  | 0.30      |+/-0.05 |milliJy             |3.81E+13|  3.00E-04|+/-5.00E-05|Jy|2010Natur.464..733S|uncertainty|     7.872 microns   | Broad-band measurement|21 35 11.6 -01 02 52.0 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
15|8.0 microns (IRAC)  | 3.5876E+02|+/-6.1994E+00|microJy             |3.81E+13|  3.59E-04|+/-6.20E-06|Jy|2013SSTSLC4.2....0C|uncertainty|7.872      microns   | Broad-band measurement|| Flux in fixed aperture|5.8" aperture                           |From new raw data
16|8.0 microns (IRAC)  | 2.9946E+02|+/-4.7438E+00|microJy             |3.81E+13|  2.99E-04|+/-4.74E-06|Jy|2013SSTSLC4.2....0C|uncertainty|7.872      microns   | Broad-band measurement|| Flux in fixed aperture|3.8" aperture                           |From new raw data
17|24 microns (MIPS)   | 2.6       |+/-0.2  |milliJy             |1.27E+13|  2.60E-03|+/-2.00E-04|Jy|2010Natur.464..733S|uncertainty|     23.68 microns   | Broad-band measurement|21 35 11.6 -01 02 52.0 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
18|24 microns (MIPS)   | 3.4048E+03|+/-2.3743E+01|microJy             |1.27E+13|  3.40E-03|+/-2.37E-05|Jy|2013SSTSLC4.2....0C|uncertainty|23.68      microns   | Broad-band measurement|| Modelled datum|PSF fit                                 |From new raw data
19|24 microns (MIPS)   | 3.2897E+03|+/-2.0554E+01|microJy             |1.27E+13|  3.29E-03|+/-2.06E-05|Jy|2013SSTSLC4.2....0C|uncertainty|23.68      microns   | Broad-band measurement|| Flux in fixed aperture|14.7" aperture                          |From new raw data
20|70 microns (MIPS)   | 6.0       |+/-2.6  |milliJy             |4.20E+12|  6.00E-03|+/-2.60E-03|Jy|2010Natur.464..733S|uncertainty|     71.42 microns   | Broad-band measurement|21 35 11.6 -01 02 52.0 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
22|250 microns Herschel| 366       |+/-55   |milliJy             |1.20E+12|  3.66E-01|+/-5.50E-02|Jy|2010A&A...518L..35I|uncertainty|       250 microns   | Broad-band measurement|| Flux integrated from map|                                        |From new raw data
26|350 microns Herschel| 429       |+/-64   |milliJy             |8.57E+11|  4.29E-01|+/-6.40E-02|Jy|2010A&A...518L..35I|uncertainty|       350 microns   | Broad-band measurement|| Flux integrated from map|                                        |From new raw data
27|352 microns (APEX)  | 530       |+/-60   |milliJy             |8.52E+11|  5.30E-01|+/-6.00E-02|Jy|2010Natur.464..733S|uncertainty|       352 microns   | Broad-band measurement|21 35 11.6 -01 02 52.0 (J2000)| Flux in fixed aperture|                                        |From new raw data
33|434 microns (SMA)   | 430       |+/-80   |milliJy             |6.91E+11|  4.30E-01|+/-8.00E-02|Jy|2010Natur.464..733S|uncertainty|       434 microns   | Broad-band measurement|21 35 11.6 -01 02 52.0 (J2000)| Flux in fixed aperture|                                        |From new raw data
34|450 microns (SCUBA) | 480       |+/-54   |milliJy             |6.66E+11|  4.80E-01|+/-5.40E-02|Jy|2010A&A...518L..35I|uncertainty|       450 microns   | Broad-band measurement|| Flux integrated from map|                                        |From new raw data
35|500 microns Herschel| 325       |+/-49   |milliJy             |6.00E+11|  3.25E-01|+/-4.90E-02|Jy|2010A&A...518L..35I|uncertainty|       500 microns   | Broad-band measurement|| Flux integrated from map|                                        |From new raw data
45|850 microns (SCUBA) | 115       |+/-13   |milliJy             |3.53E+11|  1.15E-01|+/-1.30E-02|Jy|2010A&A...518L..35I|uncertainty|       850 microns   | Broad-band measurement|| Flux integrated from map|                                        |From new raw data
47|870 microns (APEX)  | 106.0     |+/-7.0  |milliJy             |3.45E+11|  1.06E-01|+/-7.00E-03|Jy|2010Natur.464..733S|uncertainty|       870 microns   | Broad-band measurement|21 35 11.6 -01 02 52.0 (J2000)| Flux in fixed aperture|                                        |From new raw data
55|1.2 mm (SMA)        | 25.5      |+/-4.0  |milliJy             |2.50E+11|  2.55E-02|+/-4.00E-03|Jy|2010Natur.464..733S|uncertainty|       1.2 microns   | Broad-band measurement|21 35 11.6 -01 02 52.0 (J2000)| Flux in fixed aperture|                                        |From new raw data
60|2.8 mm (PdBI)       | 1.4       |+/-0.3  |milliJy             |1.07E+11|  1.40E-03|+/-3.00E-04|Jy|2010Natur.464..733S|uncertainty|       2.8 microns   | Broad-band measurement|21 35 11.6 -01 02 52.0 (J2000)| Flux in fixed aperture|                                        |From new raw data
65|8.6 mm (GBT)        | 0.13      |+/-0.04 |milliJy             |3.49E+10|  1.30E-04|+/-4.00E-05|Jy|2010Natur.464..733S|uncertainty|       8.6 microns   | Broad-band measurement|21 35 11.6 -01 02 52.0 (J2000)| Flux in fixed aperture|                                        |From new raw data
66|3.55 cm (VLA)       | 0.240     |+/-0.030|milliJy             |8.44E+09|  2.40E-04|+/-3.00E-05|Jy|2010A&A...518L..35I|uncertainty|      3.55 cm        | Broad-band measurement|| Flux integrated from map|                                        |From new raw data
67|4.49 cm (VLA)       | 0.240     |+/-0.055|milliJy             |6.68E+09|  2.40E-04|+/-5.50E-05|Jy|2010A&A...518L..35I|uncertainty|      4.49 cm        | Broad-band measurement|| Flux integrated from map|                                        |From new raw data
