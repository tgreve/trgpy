
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-04-05T08:15:36PDT



Photometric Data for SDSS J163655.77+405910.0

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|24 microns (MIPS)   |           |<225.    |mJy             |1.27E+13|  |225.E-03|Jy|2009ApJ...694.1517D|3sigma uncertainty|     23.68 microns   | Broad-band measurement|12 37 11.89 +62 22 11.8 (J2000)| Flux integrated from map|                                        |From new raw data
2|350 microns (SPIRE) | 13.7      |+/-6.9  |mJy             |8.565e+11|13.7E-03|+/-6.9e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
3|850 microns (SCUBA) |           |<3.3    |mJy             |3.53E+11|  |3.3E-03|Jy|2005MNRAS.358..149P|3rms uncertainty|     850   microns   | Broad-band measurement|12 37 11.7 +62 22 12 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
4|1.4 GHz (VLA)       | 63        |+/-21   | microJy        |1.40E+09| 63.0E-06|+/-21.0E-06|Jy|2006MNRAS.371..963B|1 sigma|       1.4 GHz       | Broad-band measurement|16 36 55.767 +40 59 09.97 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
5|1.4 GHz (VLA)       | 48.7      |+/-4.3  | microJy        |1.40E+09| 48.7E-06|+/-4.3E-06|Jy|2006MNRAS.371..963B|1 sigma|       1.4 GHz       | Broad-band measurement|16 36 55.767 +40 59 09.97 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
