
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-06-17T16:40:18PDT



Photometric Data for BzK 21000

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|R (Keck II) AB      | 23.77     || mag                |4.62E+14|  1.13E-06||Jy|2004AJ....127.3121W|no uncertainty reported|   648.7   A         | Broad-band measurement|12 37 10.744 +62 22 34.33 (J2000)| Total flux|                                        |From new raw data
2|3.6 microns (IRAC)  | 40.00     |+/-2.00 |microJy             |8.44E+13|  4.00E-05|+/-2.00E-06|Jy|2011AJ....141....1T|rms uncertainty|     3.550 microns   | Broad-band measurement|189.294266 62.376274 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
3|4.5 microns (IRAC)  | 47.50     |+/-2.38 |microJy             |6.67E+13|  4.75E-05|+/-2.38E-06|Jy|2011AJ....141....1T|rms uncertainty|     4.493 microns   | Broad-band measurement|189.294266 62.376274 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
4|5.8 microns (IRAC)  | 39.60     |+/-2.11 |microJy             |5.23E+13|  3.96E-05|+/-2.11E-06|Jy|2011AJ....141....1T|rms uncertainty|     5.731 microns   | Broad-band measurement|189.294266 62.376274 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
5|8.0 microns (IRAC)  | 44.20     |+/-2.30 |microJy             |3.81E+13|  4.42E-05|+/-2.30E-06|Jy|2011AJ....141....1T|rms uncertainty|     7.872 microns   | Broad-band measurement|189.294266 62.376274 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
6|16 microns (IRS)    | 240.4     |+/-11.5 |microJy             |1.90E+13|  2.40E-04|+/-1.15E-05|Jy|2011AJ....141....1T|rms uncertainty|      15.8 microns   | Broad-band measurement|189.294266 62.376274 (J2000)| From fitting to map|                                        |From new raw data
7|24 microns (MIPS)   | 386.0     |+/-4.9  |microJy             |1.27E+13|  3.86E-04|+/-4.90E-06|Jy|2011AJ....141....1T|rms uncertainty|     23.68 microns   | Broad-band measurement|189.294266 62.376274 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
8|24 microns (MIPS)   | 227       |+/-39   |microJy             |1.27E+13|  2.27E-04|+/-3.90E-05|Jy|2011ApJ...726...93R|uncertainty|     23.68 microns   | Broad-band measurement|12 37 10.60 +62 22 34.6 (J2000)| Not reported in paper|                                        |Averaged from previously published data
9|24 microns (MIPS)   | 392.1     |+/-5.2  |microJy             |1.27E+13|  3.92E-04|+/-5.20E-06|Jy|2011A&A...528A..35M|uncertainty|     23.68 microns   | Broad-band measurement|12 37 10.62 +62 22 34.52 (J2000)| Flux integrated from map|                                        |From new raw data
10|70 microns (MIPS)   | 3.9       |+/-0.5  | milliJy            |4.20E+12|  3.90E-03|+/-5.00E-04|Jy|2009MNRAS.399..121C|uncertainty|     71.42 microns   | Broad-band measurement|123710.60 +622234.6 (J2000)| Flux integrated from map|                                        |From reprocessed raw data
11|70 microns (MIPS)   | 5.3       |+/-0.3  |milliJy             |4.20E+12|  5.30E-03|+/-3.00E-04|Jy|2011A&A...528A..35M|uncertainty|     71.42 microns   | Broad-band measurement|12 37 10.62 +62 22 34.52 (J2000)| Flux integrated from map|                                        |From new raw data
12|100 microns (PACS)  | 8.1       |+/-0.6  |milliJy             |3.00E+12|  8.10E-03|+/-6.00E-04|Jy|2011ApJ...740L..15M|uncertainty|       100 microns   | Broad-band measurement|| From fitting to map|                                        |From reprocessed raw data
13|160 microns (PACS)  | 15.1      |+/-1.4  |milliJy             |1.87E+12|  1.51E-02|+/-1.40E-03|Jy|2011ApJ...740L..15M|uncertainty|       160 microns   | Broad-band measurement|| From fitting to map|                                        |From reprocessed raw data
14|250 microns (SPIRE) | 23.59     |+/-1.07 |milliJy             |1.20E+12|  2.36E-02|+/-1.07E-03|Jy|2010MNRAS.409...22M|uncertainty|       250 microns   | Broad-band measurement|189.294242 62.376245 (J2000)| Flux in fixed aperture|                                        |From new raw data
15|250 microns (SPIRE) | 24.4      |+/-1.5  |milliJy             |1.20E+12|  2.44E-02|+/-1.50E-03|Jy|2011ApJ...740L..15M|uncertainty|       250 microns   | Broad-band measurement|| From fitting to map|                                        |From reprocessed raw data
16|350 microns (SPIRE) | 12.59     |+/-2.05 |milliJy             |8.57E+11|  1.26E-02|+/-2.05E-03|Jy|2010MNRAS.409...22M|uncertainty|       350 microns   | Broad-band measurement|189.294242 62.376245 (J2000)| Flux in fixed aperture|                                        |From new raw data
17|350 microns (SPIRE) | 20.1      |+/-4.7  |milliJy             |8.57E+11|  2.01E-02|+/-4.70E-03|Jy|2011ApJ...740L..15M|uncertainty|       350 microns   | Broad-band measurement|| From fitting to map|                                        |From reprocessed raw data
18|500 microns (SPIRE) | 11.6      |+/-7.4  |milliJy             |6.00E+11|  1.16E-02|+/-7.40E-03|Jy|2011ApJ...740L..15M|uncertainty|       500 microns   | Broad-band measurement|| From fitting to map|                                        |From reprocessed raw data
19|850 microns (SCUBA) ||<1.8       | milliJy            |3.53E+11||1.80E-03|Jy|2009MNRAS.399..121C|2 sigma|       850 microns   | Broad-band measurement|123710.60 +622234.6 (J2000)| Flux integrated from map|                                        |From new raw data
20|CO(2-1) (IRAM)      | 0.85      |+/-0.10 | Jy km/s            |2.31E+11|  2.59E+05|+/-3.05E+04|Jy-Hz|2008ApJ...673L..21D|uncertainty|   230.539 GHz       | Line measurement; flux integrated over line; lines measured in emission|12 37 10.60 +62 22 34.6 (J2000)| Flux integrated from map|                                        |From new raw data
21|CO[2-1] (IRAM)      | 0.64      ||Jy km/s             |2.31E+11|  1.95E+05||Jy-Hz|2010ApJ...713..686D|no uncertainty reported|   230.538 GHz       | Line measurement; flux integrated over line; lines measured in emission|12 37 10.597 +62 22 34.60 (J2000)| Flux integrated from map|                                        |From new raw data
22|CO(1-0) (VLA)       | 0.13      |+/-0.03 |Jy km/s             |1.15E+11|  1.98E+04|+/-4.57E+03|Jy-Hz|2010ApJ...718..177A|uncertainty|   115.271 GHz       | Line measurement; flux integrated over line; lines measured in emission|12 37 20.597 +62 22 34.60 (J2000)| Flux integrated from map|                                        |From new raw data
23|1.4 GHz (MERLIN)    | 38.3      |+/-10.1 | microJy            |1.40E+09|  3.83E-05|+/-1.01E-05|Jy|2009MNRAS.399..121C|uncertainty|       1.4 GHz       | Broad-band measurement|123710.60 +622234.6 (J2000)| Flux integrated from map|                                        |From new raw data
24|1.4 GHz (VLA)       | 42.8      |+/-6.7  |microJy             |1.40E+09|  4.28E-05|+/-6.70E-06|Jy|2010ApJS..188..178M|uncertainty|       1.4 GHz       | Broad-band measurement|12 37 10.60 +62 22 34.6 (J2000)| Total flux; Beam filling or dilution corrected|Major=0.0"; Minor=0.0"; PA=0 deg        |From new raw data
