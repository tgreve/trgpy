
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-06-16T16:56:29PDT



Photometric Data for HS 1700+6416:[SSE2005] MD0103

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|U_n (WHT) AB        | 26.18     |+/-0.32 |mag                 |8.33E+14|  1.22E-07|+/-3.58E-08|Jy|2005ApJ...626..698S|estimated error|    0.36   microns   | Broad-band measurement|17 01 00.209 64 11 55.576 (J2000)| Flux integrated from map|                                        |From new raw data; derived from a flux in a different bandand a color
2|G (WHT) AB          | 24.69     |+/-0.17 |mag                 |6.38E+14|  4.83E-07|+/-7.40E-08|Jy|2005ApJ...626..698S|estimated error|    0.47   microns   | Broad-band measurement|17 01 00.209 64 11 55.576 (J2000)| Flux integrated from map|                                        |From new raw data; derived from a flux in a different bandand a color
3|G (WHT)             | 24.69     ||mag                 |6.38E+14|  4.83E-07||Jy|2006ApJ...647..128E|no uncertainty reported|    0.47   microns   | Broad-band measurement|| Flux in fixed aperture|                                        |Averaged from previously published data
4|H{alpha} (Keck II)  | 4.1E-17   |+/-0.8E-17|erg s^-1^ cm^-2^    |4.57E+14|  4.10E+06|+/-8.00E+05|Jy-Hz|2006ApJ...646..107E|uncertainty|    6563   A         | Line measurement; flux integrated over line; lines measured in emission|17 01 00.21 +64 11 55.58 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
5|R (WHT) AB          | 24.23     |+/-0.14 |mag                 |4.41E+14|  7.38E-07|+/-9.51E-08|Jy|2005ApJ...626..698S|estimated error|    0.68   microns   | Broad-band measurement|17 01 00.209 64 11 55.576 (J2000)| Flux integrated from map|                                        |From new raw data
6|J (Hale/WIRC)       | 21.90     ||mag                 |2.40E+14|  2.71E-06||Jy|2006ApJ...646..107E|no uncertainty reported|    1.25   microns   | Broad-band measurement|17 01 00.21 +64 11 55.58 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data; derived from aflux in a different band and a color
7|K_s (Hale/WIRC)     | 19.94     ||mag                 |1.39E+14|  7.08E-06||Jy|2006ApJ...646..107E|no uncertainty reported|    2.15   microns   | Broad-band measurement|17 01 00.21 +64 11 55.58 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data
8|K_s (P200) AB       | 22.08     |+/-0.18 |mag                 |1.39E+14|  5.34E-06|+/-9.08E-07|Jy|2005ApJ...626..698S|estimated error|    2.15   microns   | Broad-band measurement|17 01 00.209 64 11 55.576 (J2000)| Flux integrated from map|                                        |From new raw data; derived from a flux in a different bandand a color
9|3.6 microns IRAC AB | 21.32     |+/-0.10 |mag                 |8.33E+13|  1.08E-05|+/-9.91E-07|Jy|2005ApJ...626..698S|estimated error|     3.6   microns   | Broad-band measurement|17 01 00.209 64 11 55.576 (J2000)| Flux integrated from map|                                        |From new raw data
10|4.5 microns IRAC AB | 21.23     |+/-0.10 |mag                 |6.66E+13|  1.17E-05|+/-1.08E-06|Jy|2005ApJ...626..698S|estimated error|     4.5   microns   | Broad-band measurement|17 01 00.209 64 11 55.576 (J2000)| Flux integrated from map|                                        |From new raw data
11|5.8 microns IRAC AB | 21.34     |+/-0.14 |mag                 |5.17E+13|  1.06E-05|+/-1.36E-06|Jy|2005ApJ...626..698S|estimated error|     5.8   microns   | Broad-band measurement|17 01 00.209 64 11 55.576 (J2000)| Flux integrated from map|                                        |From new raw data
