

Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2010-09-03T10:19:38PDT



Photometric Data for SMM J163554.2+661225

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|F435W (HST) AB      |  27.03   |+/-0.04|mag           |6.92E+14|  5.60e-08|+/-2.06e-09|Jy|2011ApJ...734..121S|uncertainty|      4333 A         | Broad-band measurement|189.121506 62.179565 (J2000)| Total flux|                                        |From reprocessed raw data
1|F555W (HST) AB      |  26.51   |+/-0.03|mag           |5.63E+14|  9.04e-08|+/-2.50e-09|Jy|2011ApJ...734..121S|uncertainty|      4333 A         | Broad-band measurement|189.121506 62.179565 (J2000)| Total flux|                                        |From reprocessed raw data
1|F625W (HST) AB      |  26.28   |+/-0.02|mag            |4.80E+14|  1.12e-07|+/-2.06e-09|Jy|2011ApJ...734..121S|uncertainty|      4333 A         | Broad-band measurement|189.121506 62.179565 (J2000)| Total flux|                                        |From reprocessed raw data
2|F850LP (HST)         |  26.10  |+/-0.07 | mag                |3.17E+14|1.32e-07|+/-8.50e-09|Jy|2008A&A...477...55H|3 sigma|      9445 A         | Broad-band measurement|14 00 57.530 +02 52 49.34 (J2000)| Flux in fixed aperture|                                        |From new raw data
3|HST F110W            | 26.01     |+/-0.08 |mag             |2.67195e+14| 1.43e-07|+/-1.06e-08|Jy |2011ApJ...728L...4H|uncertainty|     3.550 microns   | Broad-band measurement|09 03 11.6 +00 39 06 (J2000)| Flux in fixed aperture|                                        |From new raw data
6|F160W (HST/NICMOS)  | 25.03    |+/-0.02| mag                |1.87E+14| 3.53e-07 |+/-6.51e-09|Jy|2007A&A...470..467C|internal error|       1.6 microns   | Broad-band measurement| | From fitting to map|                                        |From new raw data
21|450 microns (SCUBA) | 45        |+/-9    |milliJy             |6.66E+11|  45.0E-03|+/-9.0E-03|Jy|2006MNRAS.368..487K|uncertainty|     450   microns   | Broad-band measurement|163554.2 +661225 (J2000)| Flux integrated from map|                                        |From new raw data
21|450 microns (SCUBA) | 31.8      |+/-9.5  |milliJy             |6.66E+11|  31.8E-03|+/-9.5E-03|Jy|2006MNRAS.368..487K|uncertainty|     450   microns   | Broad-band measurement|163554.2 +661225 (J2000)| Flux integrated from map|                                        |From new raw data
25|850 microns (SCUBA) | 11        |+/-1    |milliJy             |3.53E+11|  11.0E-03|+/-1.0E-03|Jy|2006MNRAS.368..487K|uncertainty|     850   microns   | Broad-band measurement|163554.2 +661225 (J2000)| Flux integrated from map|                                        |From new raw data
25|850 microns (SCUBA) | 12.5      |+/-0.8  |milliJy             |3.53E+11|  12.8E-03|+/-1.5E-03|Jy|2006MNRAS.368..487K|uncertainty|     850   microns   | Broad-band measurement|163554.2 +661225 (J2000)| Flux integrated from map|                                        |From new raw data
