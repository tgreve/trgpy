
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-06-17T16:51:33PDT



Photometric Data for NVSS J012142+132058

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|N V 1240 (VLT)      ||<0.094E-16 |erg/s/cm^2^         |2.42E+15||9.40E+05|Jy-Hz|2009A&A...503..721M|3 sigma|      1240 A         | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|                                        |From new raw data; Extinction-corrected for Milky Way
2|C IV 1549 (VLT)     | 0.263E-16 |+/-0.005E-16|erg/s/cm^2^         |1.94E+15|  2.63E+06|+/-5.00E+04|Jy-Hz|2009A&A...503..721M|estimated error|      1549 A         | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|                                        |From new raw data; Extinction-corrected for Milky Way
3|He II 1640 (VLT)    | 0.330E-16 |+/-0.012E-16|erg/s/cm^2^         |1.83E+15|  3.30E+06|+/-1.20E+05|Jy-Hz|2009A&A...503..721M|estimated error|      1640 A         | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|                                        |From new raw data; Extinction-corrected for Milky Way
4|C III] 1909 (VLT)   | 0.282E-16 |+/-0.009E-16|erg/s/cm^2^         |1.57E+15|  2.82E+06|+/-9.00E+04|Jy-Hz|2009A&A...503..721M|estimated error|      1909 A         | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|                                        |From new raw data; Extinction-corrected for Milky Way
5|H{beta} (VLT)       | 1.0E-17   || erg/s/cm^2^        |6.17E+14|  1.00E+06||Jy-Hz|2007A&A...475..145N|no uncertainty reported|      4861 A         | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|Eastern emission line region            |From new raw data
6|H{beta} (VLT)       | 0.3E-17   || erg/s/cm^2^        |6.17E+14|  3.00E+05||Jy-Hz|2007A&A...475..145N|no uncertainty reported|      4861 A         | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|Western emission line region            |From new raw data
7|[O III] 5007 (VLT)  | 13.2E-17  || erg/s/cm^2^        |5.99E+14|  1.32E+07||Jy-Hz|2007A&A...475..145N|no uncertainty reported|      5007 A         | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|Eastern emission line region            |From new raw data
8|[O III] 5007 (VLT)  | 2.4E-17   || erg/s/cm^2^        |5.99E+14|  2.40E+06||Jy-Hz|2007A&A...475..145N|no uncertainty reported|      5007 A         | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|Western emission line region            |From new raw data
9|3.6 microns (IRAC)  | 10.5      |+/-1.8  | microJy            |8.44E+13|  1.05E-05|+/-1.80E-06|Jy|2007ApJS..171..353S|uncertainty|   3.550   microns   | Broad-band measurement|01 21 42.7 +13 20 58.00 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
10|4.5 microns (IRAC)  | 14.4      |+/-2.1  | microJy            |6.67E+13|  1.44E-05|+/-2.10E-06|Jy|2007ApJS..171..353S|uncertainty|   4.493   microns   | Broad-band measurement|01 21 42.7 +13 20 58.00 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
11|5.8 microns (IRAC)  ||<32.5      | microJy            |5.23E+13||3.25E-05|Jy|2007ApJS..171..353S|3 sigma|   5.731   microns   | Broad-band measurement|01 21 42.7 +13 20 58.00 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
12|8.0 microns (IRAC)  ||<40.3      | microJy            |3.81E+13||4.03E-05|Jy|2007ApJS..171..353S|3 sigma|   7.872   microns   | Broad-band measurement|01 21 42.7 +13 20 58.00 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
13|16 microns (IRS)    ||<136.0     | microJy            |1.87E+13||1.36E-04|Jy|2007ApJS..171..353S|3 sigma|      16   microns   | Broad-band measurement|01 21 42.7 +13 20 58.00 (J2000)| Flux in fixed aperture|6" diameter aperture                    |From reprocessed raw data
14|450 microns (SCUBA) | 4         |+/-16   | milliJy            |6.66E+11|  4.00E-03|+/-1.60E-02|Jy|2004MNRAS.353..377R|uncertainty|       450 microns   | Broad-band measurement|01 21 42.74 +13 20 58.3 (J2000)| Not reported in paper|Good quality data                       |From new raw data
15|850 microns (SCUBA) | 7.5       |+/-1.0  |milliJy             |3.53E+11|  7.50E-03|+/-1.00E-03|Jy|2007MNRAS.375.1299V|uncertainty|     850   microns   | Broad-band measurement|| Flux integrated from map|From 2001MNRAS.323..417A                |Averaged from previously published data
16|850 microns (SCUBA) | 7.5       |+/-1.0  | milliJy            |3.53E+11|  7.50E-03|+/-1.00E-03|Jy|2004MNRAS.353..377R|uncertainty|       850 microns   | Broad-band measurement|01 21 42.74 +13 20 58.3 (J2000)| Not reported in paper|Good quality data                       |From new raw data
17|1.4GHz              | 55.4      |+/-1.7  |milliJy             |1.40E+09|  5.54E-02|+/-1.70E-03|Jy|1998AJ....115.1693C|uncertainty|    1.40   GHz       | Broad-band measurement|01 21 42.73 +13 20 58.1 (J2000)| Flux integrated from map|                                        |From new raw data
18|365 MHz (Texas)     | 0.348     |+/-0.027|Jy                  |3.65E+08|  3.48E-01|+/-2.70E-02|Jy|1996AJ....111.1945D|internal error|365        MHz       | Broad-band measurement; obtained by interpolation over frequency|011903.546 130516.91 (B1950)| Integrated from scans|Model:P;MFlag:+;EFlag:+;LFlag:+.        |From new raw data
19|74 MHz (VLA)        | 2.02      |+/-0.22 | Jy                 |7.38E+07|  2.02E+00|+/-2.20E-01|Jy|2007AJ....134.1245C|rms uncertainty|    73.8   MHz       | Broad-band measurement|01 21 42.60 +13 21 00.5 (J2000)| Flux integrated from map|Corrected for clean bias                |From new raw data
