
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2017-01-03T06:04:38PST



Photometric Data for SDSS J1148+5251

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|3000 A              | 4.22E-17  |+/-0.08E-17|erg/s/cm^2^/A       |9.99E+14|  1.27E-05|+/-2.41E-07|Jy|2011ApJ...739...56D|uncertainty|      3000 A         | Broad-band measurement|| Modelled datum|                                        |Transformed from previously published data
2|R (Keck /LRIS) AB  | 25.2      |+/-0.3  |mag                 |4.67E+14|  3.02E-07|+/-8.35E-08|Jy|2005ApJ...634L...9M|estimated error|    6417   A         | Broad-band measurement|11 48 16.67 +52 51 50.4 (J2000)| Flux in fixed aperture|2.5" diameter aperture                  |From new raw data
3|i (PAN-STARRS1) AB  ||>23.07     |mag                 |3.97E+14||2.15E-06|Jy|2014AJ....148...14B|3 sigma|      7549 A         | Broad-band measurement|11 48 16.65 +52 51 50.4 (J2000)| Flux in fixed aperture|                                        |From new raw data
4|F775W (HST/ACS) AB      | 22.86     ||mag                 |3.86E+14|  2.61E-06||Jy|2009ApJ...695..809K|no uncertainty reported|      7764 A         | Broad-band measurement|11 48 16.74 +52 51 50.11 (J2000)| Flux in fixed aperture|                                        |From new raw data; derived from a flux in a different bandand a color
5|z (PAN-STARRS1) AB  | 20.63     |+/-0.04 |mag                 |3.45E+14|  2.03E-05|+/-7.49E-07|Jy|2014AJ....148...14B|uncertainty|      8701 A         | Broad-band measurement|11 48 16.65 +52 51 50.4 (J2000)| Flux in fixed aperture|                                        |From new raw data
6|z (Keck /LRIS) AB  | 19.7      |+/-0.3  |mag                 |3.30E+14|  4.79E-05|+/-1.32E-05|Jy|2005ApJ...634L...9M|estimated error|    9097   A         | Broad-band measurement|11 48 16.67 +52 51 50.4 (J2000)| Flux in fixed aperture|2.5" diameter aperture                  |From new raw data
7|F850LP (HST/ACS) AB     | 19.83     ||mag                 |3.17E+14|  4.25E-05||Jy|2009ApJ...695..809K|no uncertainty reported|      9445 A         | Broad-band measurement|11 48 16.74 +52 51 50.11 (J2000)| Total flux|                                        |From new raw data
8|y (PAN-STARRS1) AB  | 19.42     |+/-0.10 |mag                 |3.15E+14|  6.20E-05|+/-5.71E-06|Jy|2014AJ....148...14B|uncertainty|      9510 A         | Broad-band measurement|11 48 16.65 +52 51 50.4 (J2000)| Flux in fixed aperture|                                        |From new raw data
9|J (Hale/WIRC)       | 18.07     |+/-0.02 |mag                 |2.40E+14|  9.42E-05|+/-1.73E-06|Jy|2005ApJ...634L...9M|uncertainty|    1.25   microns   | Broad-band measurement|11 48 16.67 +52 51 50.4 (J2000)| Flux in fixed aperture|3.5" diameter aperture                  |From new raw data
10|H (Subaru)          | 17.70     |+/-0.05 |mag                 |1.83E+14|  8.48E-05|+/-3.91E-06|Jy|2004ApJ...614...69I|typical accuracy|      1.64 microns   | Broad-band measurement|114816.64 +525150.3 (J2000)| Flux in fixed aperture|2.2" diameter aperture                  |From new raw data
11|K' (Subaru)         | 16.98     |+/-0.05 |mag                 |1.41E+14|  1.15E-04|+/-5.28E-06|Jy|2004ApJ...614...69I|typical accuracy|      2.13 microns   | Broad-band measurement|114816.64 +525150.3 (J2000)| Flux in fixed aperture|2.2" diameter aperture                  |From new raw data
12|K (Keck)            | 18.1      || mag                |1.37E+14|  3.57E-05||Jy|2009MNRAS.395.1476R|no uncertainty reported|      2.19 microns   | Broad-band measurement|| Not reported in paper|                                        |From new raw data
13|3.6 microns (IRAC)  | 1.0971E+02|+/-1.4688E-01|microJy             |8.44E+13|  1.10E-04|+/-1.47E-07|Jy|2013SSTSLC4.2....0C|uncertainty|3.55       microns   | Broad-band measurement|| Flux in fixed aperture|3.8" aperture                           |From new raw data
14|3.6 microns (IRAC)  | 1.3082E+02|+/-2.9199E-01|microJy             |8.44E+13|  1.31E-04|+/-2.92E-07|Jy|2013SSTSLC4.2....0C|uncertainty|3.55       microns   | Broad-band measurement|| Flux in fixed aperture|3.8" aperture                           |From new raw data
15|3.6 microns (IRAC)  | 1.2885E+02|+/-3.4200E-01|microJy             |8.44E+13|  1.29E-04|+/-3.42E-07|Jy|2013SSTSLC4.2....0C|uncertainty|3.55       microns   | Broad-band measurement|| Flux in fixed aperture|5.8" aperture                           |From new raw data
16|3.6 microns (IRAC)  | 1.3237E+02|+/-2.5434E-01|microJy             |8.44E+13|  1.32E-04|+/-2.54E-07|Jy|2013SSTSLC4.2....0C|uncertainty|3.55       microns   | Broad-band measurement|| Flux in fixed aperture|5.8" aperture                           |From new raw data
17|3.6 microns (IRAC)  | 0.124     |+/-0.002|milliJy             |8.44E+13|  1.24E-04|+/-2.00E-06|Jy|2006AJ....132.2127J|uncertainty|   3.550   microns   | Broad-band measurement|| Flux in fixed aperture|6 pixel aper; bkgd annulus 8-13 pixels  |From reprocessed raw data
18|4.5 microns (IRAC)  | 1.4970E+02|+/-5.1187E-01|microJy             |6.67E+13|  1.50E-04|+/-5.12E-07|Jy|2013SSTSLC4.2....0C|uncertainty|4.493      microns   | Broad-band measurement|| Flux in fixed aperture|5.8" aperture                           |From new raw data
19|4.5 microns (IRAC)  | 1.1009E+02|+/-3.9028E-01|microJy             |6.67E+13|  1.10E-04|+/-3.90E-07|Jy|2013SSTSLC4.2....0C|uncertainty|4.493      microns   | Broad-band measurement|| Flux in fixed aperture|3.8" aperture                           |From new raw data
20|4.5 microns (IRAC)  | 1.4392E+02|+/-2.8315E-01|microJy             |6.67E+13|  1.44E-04|+/-2.83E-07|Jy|2013SSTSLC4.2....0C|uncertainty|4.493      microns   | Broad-band measurement|| Flux in fixed aperture|3.8" aperture                           |From new raw data
21|4.5 microns (IRAC)  | 1.2124E+02|+/-5.7253E-01|microJy             |6.67E+13|  1.21E-04|+/-5.73E-07|Jy|2013SSTSLC4.2....0C|uncertainty|4.493      microns   | Broad-band measurement|| Flux in fixed aperture|5.8" aperture                           |From new raw data
22|4.5 microns (IRAC)  | 0.140     |+/-0.003|milliJy             |6.67E+13|  1.40E-04|+/-3.00E-06|Jy|2006AJ....132.2127J|uncertainty|   4.493   microns   | Broad-band measurement|| Flux in fixed aperture|6 pixel aper; bkgd annulus 8-13 pixels  |From reprocessed raw data
23|5.8 microns (IRAC)  | 1.3807E+02|+/-1.9914E+00|microJy             |5.23E+13|  1.38E-04|+/-1.99E-06|Jy|2013SSTSLC4.2....0C|uncertainty|5.731      microns   | Broad-band measurement|| Flux in fixed aperture|5.8" aperture                           |From new raw data
24|5.8 microns (IRAC)  | 1.2088E+02|+/-1.3383E+00|microJy             |5.23E+13|  1.21E-04|+/-1.34E-06|Jy|2013SSTSLC4.2....0C|uncertainty|5.731      microns   | Broad-band measurement|| Flux in fixed aperture|3.8" aperture                           |From new raw data
25|5.8 microns (IRAC)  | 1.3903E+02|+/-2.1020E+00|microJy             |5.23E+13|  1.39E-04|+/-2.10E-06|Jy|2013SSTSLC4.2....0C|uncertainty|5.731      microns   | Broad-band measurement|| Flux in fixed aperture|5.8" aperture                           |From new raw data
26|5.8 microns (IRAC)  | 1.4355E+02|+/-1.5327E+00|microJy             |5.23E+13|  1.44E-04|+/-1.53E-06|Jy|2013SSTSLC4.2....0C|uncertainty|5.731      microns   | Broad-band measurement|| Flux in fixed aperture|3.8" aperture                           |From new raw data
27|5.8 microns (IRAC)  | 0.133     |+/-0.010|milliJy             |5.23E+13|  1.33E-04|+/-1.00E-05|Jy|2006AJ....132.2127J|uncertainty|   5.731   microns   | Broad-band measurement|| Flux in fixed aperture|6 pixel aper; bkgd annulus 8-13 pixels  |From reprocessed raw data
28|8.0 microns (IRAC)  | 0.241     |+/-0.016|milliJy             |3.81E+13|  2.41E-04|+/-1.60E-05|Jy|2006AJ....132.2127J|uncertainty|   7.872   microns   | Broad-band measurement|| Flux in fixed aperture|6 pixel aper; bkgd annulus 8-13 pixels  |From reprocessed raw data
29|8.0 microns (IRAC)  | 2.0452E+02|+/-3.1410E+00|microJy             |3.81E+13|  2.05E-04|+/-3.14E-06|Jy|2013SSTSLC4.2....0C|uncertainty|7.872      microns   | Broad-band measurement|| Flux in fixed aperture|5.8" aperture                           |From new raw data
30|8.0 microns (IRAC)  | 1.9218E+02|+/-3.0397E+00|microJy             |3.81E+13|  1.92E-04|+/-3.04E-06|Jy|2013SSTSLC4.2....0C|uncertainty|7.872      microns   | Broad-band measurement|| Flux in fixed aperture|5.8" aperture                           |From new raw data
31|8.0 microns (IRAC)  | 1.7220E+02|+/-2.2110E+00|microJy             |3.81E+13|  1.72E-04|+/-2.21E-06|Jy|2013SSTSLC4.2....0C|uncertainty|7.872      microns   | Broad-band measurement|| Flux in fixed aperture|3.8" aperture                           |From new raw data
32|8.0 microns (IRAC)  | 2.0837E+02|+/-2.3887E+00|microJy             |3.81E+13|  2.08E-04|+/-2.39E-06|Jy|2013SSTSLC4.2....0C|uncertainty|7.872      microns   | Broad-band measurement|| Flux in fixed aperture|3.8" aperture                           |From new raw data
33|16 microns (IRS/Spitzer)| 0.51      |+/-10  %| milliJy            |1.86E+13|  5.10E-04|+/-5.10E-05|Jy|2004ApJS..154..142C|uncertainty|     16.10 microns   | Broad-band measurement|11 48 16.5 +52 51 49.1 (J2000)| Flux integrated from map|                                        |From new raw data
34|22 microns (IRS/Spitzer)| 0.74      |+/-10  %| milliJy            |1.35E+13|  7.40E-04|+/-7.40E-05|Jy|2004ApJS..154..142C|uncertainty|     22.25 microns   | Broad-band measurement|11 48 16.5 +52 51 49.1 (J2000)| Flux integrated from map|                                        |From new raw data
35|24 microns (MIPS)   | 1.520     |+/-0.130|milliJy             |1.27E+13|  1.52E-03|+/-1.30E-04|Jy|2006AJ....132.2127J|uncertainty|   23.68   microns   | Broad-band measurement|| Flux in fixed aperture|6 pixel aper; bkgd annulus 8-13 pixels  |Averaged from previously published data
36|24 microns (MIPS)   | 1.52      |+/-0.12 |milliJy             |1.27E+13|  1.52E-03|+/-1.20E-04|Jy|2006ApJ...641L..85H|estimated error|   23.68   microns   | Broad-band measurement|| Corrected to total flux from single aperture measurement|Absolute calibration uncertainty is 10% |From new raw data
37|24 microns (MIPS)   | 1.3343E+03|+/-2.5033E+01|microJy             |1.27E+13|  1.33E-03|+/-2.50E-05|Jy|2013SSTSLC4.2....0C|uncertainty|23.68      microns   | Broad-band measurement|| Modelled datum|PSF fit                                 |From new raw data
38|24 microns (MIPS)   | 1.2735E+03|+/-2.3002E+01|microJy             |1.27E+13|  1.27E-03|+/-2.30E-05|Jy|2013SSTSLC4.2....0C|uncertainty|23.68      microns   | Broad-band measurement|| Flux in fixed aperture|14.7" aperture                          |From new raw data
39|70 microns (MIPS)   ||<9.73      |milliJy             |4.20E+12||9.73E-03|Jy|2006AJ....132.2127J|2 sigma|   71.42   microns   | Broad-band measurement|| Flux in fixed aperture|35" aperture; 39"-65" bkgd annulus      |From reprocessed raw data
40|100 microns (PACS)  | 4.1       |+/-1.0  |milliJy             |3.00E+12|  4.10E-03|+/-1.00E-03|Jy|2010A&A...518L..34L|uncertainty|     100.0 microns   | Broad-band measurement|| Flux in fixed aperture|5.0" radius aperture                    |From new raw data
41|160 microns (PACS)  | 6.3       |+/-2.0  |milliJy             |1.87E+12|  6.30E-03|+/-2.00E-03|Jy|2010A&A...518L..34L|uncertainty|     160.0 microns   | Broad-band measurement|| Flux in fixed aperture|5.0" radius aperture                    |From new raw data
42|[N II] (IRAM)       ||<0.48      | Jy km/s            |1.46E+12||3.15E+05|Jy-Hz|2009ApJ...691L...1W|3 sigma|  1461.132 GHz       | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|                                        |From new raw data
43|350 microns SHARC II| 21        |+/-6    |milliJy             |8.57E+11|  2.10E-02|+/-6.00E-03|Jy|2006ApJ...642..694B|1 sigma|     350   microns   | Broad-band measurement|11 48 16.64 +52 51 50.30 (J2000)| Flux integrated from map|                                        |From new raw data
44|CO(7-6) (PdBI)      | 0.63      |+/-0.06 |Jy km/s             |8.07E+11|  2.29E+05|+/-2.18E+04|Jy-Hz|2009ApJ...703.1338R|uncertainty|    806.65 GHz       | Line measurement; flux integrated over line; lines measured in emission|11 48 16.64 +52 51 50.3 (J2000)| Flux integrated from map|                                        |From new raw data
45|CO(6-5) (IRAM)      | 1.12      |+/-0.3  | Jy km/s            |6.91E+11|  3.48E+05|+/-9.33E+04|Jy-Hz|2009ApJ...691L...1W|uncertainty|   691.473 GHz       | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|                                        |From new raw data
46|450 microns (SCUBA) | 24.7      |+/-7.4  |milliJy             |6.66E+11|  2.47E-02|+/-7.40E-03|Jy|2004MNRAS.351L..29R|1 sigma|     450   microns   | Broad-band measurement|11 48 16.64 +52 51 50.3 (J2000)| Flux integrated from map|                                        |From new raw data
47|850 microns (SCUBA) | 7.8       |+/-0.7  |milliJy             |3.53E+11|  7.80E-03|+/-7.00E-04|Jy|2004MNRAS.351L..29R|1 sigma|     850   microns   | Broad-band measurement|11 48 16.64 +52 51 50.3 (J2000)| Flux integrated from map|                                        |From new raw data
48|HCN(J=2-1) (VLA)    ||<30        | microJy            |1.77E+11||3.20E-05|Jy|2007ApJ...671L..13R|2 sigma|   177.261 GHz       | Line measurement; flux integrated over line|| Peak flux|                                        |From new raw data
49|46.6 GHz (VLA)      ||<0.10      | milliJy            |4.66E+10||1.00E-04|Jy|2004ApJ...615L..17W|2 sigma|     46.61 GHz       | Broad-band measurement|| Flux integrated from map|From 2003Natur.424..406W                |Averaged from previously published data
50|23.9 GHz (VLA)      ||<22        | microJy            |2.39E+10||2.20E-05|Jy|2007ApJ...671L..13R|2 sigma|     23.89 GHz       | Broad-band measurement|| Peak flux|                                        |From new raw data
51|1.4 GHz (VLA)       | 55        |+/-12   | microJy            |1.40E+09|  5.50E-05|+/-1.20E-05|Jy|2004AJ....128..997C|uncertainty|       1.4 GHz       | Broad-band measurement|11 48 16.65 +52 51 50.2 (J2000)| Flux integrated from map|4.6 sigma detection                     |From new raw data
