\queryDateTime = 2018-11-27T11:57:07PST
\source = /hydra/workarea/irsaviewer/temp_files/IpacTableFromSource2257050731345606935.tbl
\QUERY_STATUS = OK
\CatalogTargetColName = Coordinates Targeted
\Description = Published and Homogenized [Frequency, Flux Dens...
\LINK = http://ned.ipac.caltech.edu/cgi-bin/datasearch?sea
\
z=0.00298
|No.   |Observed Passband   |Photometry Measurement|Uncertainty  |Units            |Frequency|Flux Density|Upper limit of uncertainty|Lower limit of uncertainty|Upper limit of Flux Density|Lower limit of Flux Density|NED Uncertainty|NED Units|Refcode            |Significance           |Published frequency|Frequency Mode                                                                              |Coordinates Targeted           |Spatial Mode                                            |Qualifiers                             |Comments                                                                                                                                                           |
|int   |char                |double                |char         |char             |double   |double      |double                    |double                    |double                     |double                     |char           |char     |char               |char                   |char               |char                                                                                        |char                           |char                                                    |char                                   |char                                                                                                                                                               |
|      |                    |                      |             |                 |Hz       |Jy          |                          |                          |                           |                           |               |         |                   |                       |                   |                                                                                            |                               |                                                        |                                       |                                                                                                                                                                   |
|      |                    |                      |             |                 |         |            |                          |                          |                           |                           |               |         |                   |                       |                   |                                                                                            |                               |                                                        |                                       |                                                                                                                                                                   |
 1     |2-10 keV (Chandra)  |9.8E-13               |             |erg/cm^2^/s      |1.45E+18 |6.76E-08    |                          |                          |                           |                           |               |Jy       |2005PASJ...57..135I|no uncertainty reported|6   keV            |Broad-band measurement                                                                      |                               |Total flux                                              |                                       |From new raw data; NED frequency assigned to mid-point ofband in keV                                                                                               
 2     |0.2-10 keV (Chandra)|5.5E-15               |             |ergs/cm^2^/s     |1.23E+18 |4.45E-10    |                          |                          |                           |                           |               |Jy       |2007A&A...468..129T|no uncertainty reported|5.10   keV         |Broad-band measurement                                                                      |06 18 37.6 +78 21 20 (J2000)   |Flux integrated from map                                |                                       |From reprocessed raw data; NED frequency assigned tomid-point of band in keV                                                                                       
 3     |0.2-2 keV (ROSAT)   |6.4E-13               |+/-6.8 %     |erg/s/cm^2^      |3.15E+17 |2.03E-07    |1.38E-08                  |1.38E-08                  |                           |                           |+/-1.38E-08    |Jy       |2000WGA...C...0000W|mean error             |1.3       keV      |Broad-band measurement                                                                      |061836.9 +782121. (J2000)      |Flux integrated from map                                |                                       |From reprocessed raw data; NED frequency assigned tomid-point of band in keV                                                                                       
 4     |FUV (GALEX) AB      |1.6E+01               |+/-0.01      |mag              |1.98E+15 |2.13E-03    |1.96E-05                  |1.96E-05                  |                           |                           |+/-1.96E-05    |Jy       |2007ApJS..173..185G|uncertainty            |1516 A             |Broad-band measurement                                                                      |06 18 37.7 +78 21 25.3 (J2000) |Total flux                                              |                                       |From new raw data                                                                                                                                                  
 5     |UV_1650 (m_T)       |1.2E+01               |+/-0.30      |mag              |1.82E+15 |3.52E-03    |1.12E-03                  |1.12E-03                  |                           |                           |+/-1.12E-03    |Jy       |1995A&AS..114..527R|mean error             |1650       A       |Broad-band measurement; broad-band flux derived by integration over spectrum; synthetic band|061043 782223 (B1950)          |Multiple methods                                        |                                       |Homogenized from previously published data                                                                                                                         
 6     |NUV (GALEX) AB      |1.5E+01               |+/-0.01      |mag              |1.32E+15 |4.70E-03    |4.33E-05                  |4.33E-05                  |                           |                           |+/-4.33E-05    |Jy       |2007ApJS..173..185G|uncertainty            |2267 A             |Broad-band measurement                                                                      |06 18 37.7 +78 21 25.3 (J2000) |Total flux                                              |                                       |From new raw data                                                                                                                                                  
 7     |UV_2500 (m_T)       |1.4E+01               |+/-0.46      |mag              |1.20E+15 |2.83E-03    |1.49E-03                  |1.49E-03                  |                           |                           |+/-1.49E-03    |Jy       |1995A&AS..114..527R|mean error             |2500       A       |Broad-band measurement; broad-band flux derived by integration over spectrum; synthetic band|061043 782223 (B1950)          |Multiple methods                                        |                                       |Homogenized from previously published data                                                                                                                         
 8     |UV_3150 (m_T)       |1.2E+01               |+/-0.30      |mag              |9.52E+14 |2.75E-02    |8.76E-03                  |8.76E-03                  |                           |                           |+/-8.76E-03    |Jy       |1995A&AS..114..527R|mean error             |3150       A       |Broad-band measurement; broad-band flux derived by integration over spectrum; synthetic band|061043 782223 (B1950)          |Multiple methods                                        |                                       |Homogenized from previously published data                                                                                                                         
 9     |U (U_T^0)           |1.1E+01               |             |mag              |8.19E+14 |9.07E-02    |                          |                          |                           |                           |               |Jy       |1991RC3.9.C...0000d|no uncertainty reported|3660       A       |Broad-band measurement                                                                      |061042.7 +782223 (B1950)       |From multi-aperture data                                |                                       |Homogenized from new and previously published data;Extinction-corrected for internal and Milky Way and K-correction applied; Standard Johnson UBVRI filters assumed
 10    |U (U_T)             |1.2E+01               |+/-0.14      |mag              |8.19E+14 |3.89E-02    |5.19E-03                  |5.19E-03                  |                           |                           |+/-5.19E-03    |Jy       |1991RC3.9.C...0000d|rms uncertainty        |3660       A       |Broad-band measurement                                                                      |061042.7 +782223 (B1950)       |From multi-aperture data                                |                                       |Homogenized from new and previously published data; StandardJohnson UBVRI filters assumed                                                                          
 17    |B (B_T)             |1.1E+01               |+/-0.13      |mag              |6.81E+14 |1.20E-01    |1.52E-02                  |1.52E-02                  |                           |                           |+/-1.52E-02    |Jy       |1991RC3.9.C...0000d|rms uncertainty        |4400       A       |Broad-band measurement                                                                      |061042.7 +782223 (B1950)       |From multi-aperture data                                |                                       |Homogenized from new and previously published data; StandardJohnson UBVRI filters assumed                                                                          
 18    |B (B_T^0)           |1.1E+01               |             |mag              |6.81E+14 |2.50E-01    |                          |                          |                           |                           |               |Jy       |1991RC3.9.C...0000d|no uncertainty reported|4400       A       |Broad-band measurement                                                                      |061042.7 +782223 (B1950)       |Multiple methods                                        |                                       |Homogenized from new and previously published data;Extinction-corrected for internal and Milky Way and K-correction applied; Standard Johnson UBVRI filters assumed
 19    |m_p                 |1.1E+01               |+/-0.4       |mag              |6.81E+14 |1.55E-01    |6.89E-02                  |6.89E-02                  |                           |                           |+/-6.89E-02    |Jy       |1968CGCG4.C...0000Z|rms noise              |4400       A       |Broad-band measurement                                                                      |061030.0 +782200. (B1950)      |Estimated by eye                                        |                                       |From new raw data                                                                                                                                                  
 20    |B (Cousins)         |1.1E+01               |+/-0.02      |mag              |6.81E+14 |1.16E-01    |2.16E-03                  |2.16E-03                  |                           |                           |+/-2.16E-03    |Jy       |1996A&AS..118..111H|uncertainty            |4400       A       |Broad-band measurement                                                                      |06 17 52.5 +78 21 27 (1995 )   |Flux in fixed aperture                                  |                                       |From new raw data                                                                                                                                                  
 21    |B (m_B)             |1.1E+01               |+/-0.14      |mag              |6.81E+14 |1.65E-01    |2.27E-02                  |2.27E-02                  |                           |                           |+/-2.27E-02    |Jy       |1991RC3.9.C...0000d|rms uncertainty        |4400       A       |Broad-band measurement                                                                      |061042.7 +782223 (B1950)       |Multiple methods                                        |                                       |Homogenized from new and previously published data; StandardJohnson UBVRI filters assumed                                                                          
 26    |V (Cousins)         |1.1E+01               |+/-0.06      |mag              |5.45E+14 |1.89E-01    |1.08E-02                  |1.08E-02                  |                           |                           |+/-1.08E-02    |Jy       |1996A&AS..118..111H|uncertainty            |5500       A       |Broad-band measurement                                                                      |06 17 52.5 +78 21 27 (1995 )   |Flux in fixed aperture                                  |                                       |From new raw data                                                                                                                                                  
 27    |V (Johnson)         |1.3E+01               |             |mag              |5.42E+14 |1.76E-02    |                          |                          |                           |                           |               |Jy       |1988VIrPh.C...0000d|no uncertainty reported|5530   A           |Broad-band measurement                                                                      |                               |Flux in fixed aperture                                  |25" aperture                           |Transformed from previously published data; Standard JohnsonUBVRI filters assumed                                                                                  
 28    |V (V_T^0)           |1.0E+01               |             |mag              |5.42E+14 |3.81E-01    |                          |                          |                           |                           |               |Jy       |1991RC3.9.C...0000d|no uncertainty reported|5530       A       |Broad-band measurement                                                                      |061042.7 +782223 (B1950)       |From multi-aperture data                                |                                       |Homogenized from new and previously published data;Extinction-corrected for internal and Milky Way and K-correction applied; Standard Johnson UBVRI filters assumed
 29    |V (V_T)             |1.1E+01               |+/-0.13      |mag              |5.42E+14 |2.11E-01    |2.72E-02                  |2.72E-02                  |                           |                           |+/-2.72E-02    |Jy       |1991RC3.9.C...0000d|rms uncertainty        |5530       A       |Broad-band measurement                                                                      |061042.7 +782223 (B1950)       |From multi-aperture data                                |                                       |Homogenized from new and previously published data; StandardJohnson UBVRI filters assumed                                                                          
 30    |R (Johnson) (IAC80) |9.8E+00               |+/-0.05      |mag              |5.00E+14 |3.38E-01    |1.56E-02                  |1.56E-02                  |                           |                           |+/-1.56E-02    |Jy       |2004AJ....127.1386C|uncertainty            |6000   A           |Broad-band measurement                                                                      |                               |Flux in fixed aperture                                  |159.16" circular aperture radius       |From new raw data                                                                                                                                                  
 33    |R (Johnson) (JKT)   |1.0E+01               |+/-0.04      |mag              |4.70E+14 |2.74E-01    |1.01E-02                  |1.01E-02                  |                           |                           |+/-1.01E-02    |Jy       |2004A&A...414...23J|uncertainty            |6373   A           |Broad-band measurement                                                                      |                               |Total flux                                              |                                       |From new raw data                                                                                                                                                  
 44    |R (Johnson)         |1.2E+01               |             |mag              |4.28E+14 |4.25E-02    |                          |                          |                           |                           |               |Jy       |1988VIrPh.C...0000d|no uncertainty reported|7000   A           |Broad-band measurement                                                                      |                               |Flux in fixed aperture                                  |25" aperture                           |Transformed from previously published data; Standard JohnsonUBVRI filters assumed                                                                                  
 45    |I (Cousins)         |9.6E+00               |+/-0.14      |mag              |3.79E+14 |3.55E-01    |4.89E-02                  |4.89E-02                  |                           |                           |+/-4.89E-02    |Jy       |1996A&AS..118..111H|uncertainty            |7900       A       |Broad-band measurement                                                                      |06 17 52.5 +78 21 27 (1995 )   |Flux in fixed aperture                                  |                                       |From new raw data                                                                                                                                                  
 46    |I (Johnson) (IAC80) |9.2E+00               |+/-0.06      |mag              |3.41E+14 |4.68E-01    |2.58E-02                  |2.58E-02                  |                           |                           |+/-2.58E-02    |Jy       |2004AJ....127.1386C|uncertainty            |8800   A           |Broad-band measurement                                                                      |                               |Flux in fixed aperture                                  |168.67" circular aperture radius       |From new raw data                                                                                                                                                  
 47    |J (Johnson)         |8.6E+00               |+/-0.03      |mag              |2.42E+14 |5.98E-01    |1.68E-02                  |1.68E-02                  |                           |                           |+/-1.68E-02    |Jy       |1977HarvU.T00M....A|uncertainty            |1.24    microns    |Broad-band measurement                                                                      |                               |Flux in fixed aperture                                  |105" aperture                          |From new raw data; derived from a flux in a different bandand a color                                                                                              
 48    |J (Johnson)         |9.7E+00               |+/-0.03      |mag              |2.42E+14 |2.21E-01    |6.20E-03                  |6.20E-03                  |                           |                           |+/-6.20E-03    |Jy       |1977HarvU.T00M....A|uncertainty            |1.24    microns    |Broad-band measurement                                                                      |                               |Flux in fixed aperture                                  |27.4" aperture                         |From new raw data; derived from a flux in a different bandand a color                                                                                              
 49    |J (Johnson)         |9.2E+00               |+/-0.03      |mag              |2.42E+14 |3.29E-01    |9.21E-03                  |9.21E-03                  |                           |                           |+/-9.21E-03    |Jy       |1977HarvU.T00M....A|uncertainty            |1.24    microns    |Broad-band measurement                                                                      |                               |Flux in fixed aperture                                  |41.1" aperture                         |From new raw data; derived from a flux in a different bandand a color                                                                                              
 50    |J_14arcsec (2MASS)  |1.0E+01               |+/-0.015     |mag              |2.40E+14 |1.20E-01    |1.67E-03                  |1.67E-03                  |                           |                           |+/-1.67E-03    |Jy       |20032MASX.C.......:|1 sigma uncert.        |1.25      microns  |Broad-band measurement                                                                      |061837.71 +782125.3 (J2000)    |Flux in fixed aperture                                  |14.0 x 14.0 arcsec aperture            |From new raw data                                                                                                                                                  
 51    |J_Kron (2MASS LGA)  |8.4E+00               |+/-0.015     |mag              |2.40E+14 |6.65E-01    |9.26E-03                  |9.26E-03                  |                           |                           |+/-9.26E-03    |Jy       |2003AJ....125..525J|1 sigma uncert.        |1.25      microns  |Broad-band measurement                                                                      |061837.71 +782125.3 (J2000)    |Flux integrated from map                                |174.8 x   82.2 arcsec integration area.|From new raw data; Corrected for contaminating sources                                                                                                             
 52    |J_tot (2MASS LGA)   |8.2E+00               |+/-0.020     |mag              |2.40E+14 |8.14E-01    |1.51E-02                  |1.51E-02                  |                           |                           |+/-1.51E-02    |Jy       |2003AJ....125..525J|1 sigma uncert.        |1.25      microns  |Broad-band measurement                                                                      |061837.71 +782125.3 (J2000)    |Total flux                                              |                                       |From new raw data                                                                                                                                                  
 53    |J_20 (2MASS LGA)    |8.4E+00               |+/-0.016     |mag              |2.40E+14 |6.98E-01    |1.04E-02                  |1.04E-02                  |                           |                           |+/-1.04E-02    |Jy       |2003AJ....125..525J|1 sigma uncert.        |1.25      microns  |Broad-band measurement                                                                      |061837.71 +782125.3 (J2000)    |Flux integrated from map                                |195.0 x   91.7 arcsec integration area.|From new raw data; Corrected for contaminating sources                                                                                                             
 54    |H_14arcsec (2MASS)  |9.2E+00               |+/-0.015     |mag              |1.82E+14 |2.12E-01    |2.95E-03                  |2.95E-03                  |                           |                           |+/-2.95E-03    |Jy       |20032MASX.C.......:|1 sigma uncert.        |1.65      microns  |Broad-band measurement                                                                      |061837.71 +782125.3 (J2000)    |Flux in fixed aperture                                  |14.0 x 14.0 arcsec aperture            |From new raw data                                                                                                                                                  
 55    |H_tot (2MASS LGA)   |7.4E+00               |+/-0.021     |mag              |1.82E+14 |1.11E+00    |2.16E-02                  |2.16E-02                  |                           |                           |+/-2.16E-02    |Jy       |2003AJ....125..525J|1 sigma uncert.        |1.65      microns  |Broad-band measurement                                                                      |061837.71 +782125.3 (J2000)    |Total flux                                              |                                       |From new raw data                                                                                                                                                  
 56    |H_20 (2MASS LGA)    |7.6E+00               |+/-0.016     |mag              |1.82E+14 |9.72E-01    |1.44E-02                  |1.44E-02                  |                           |                           |+/-1.44E-02    |Jy       |2003AJ....125..525J|1 sigma uncert.        |1.65      microns  |Broad-band measurement                                                                      |061837.71 +782125.3 (J2000)    |Flux integrated from map                                |195.0 x   91.7 arcsec integration area.|From new raw data; Corrected for contaminating sources                                                                                                             
 57    |H_Kron (2MASS LGA)  |7.6E+00               |+/-0.016     |mag              |1.82E+14 |9.35E-01    |1.39E-02                  |1.39E-02                  |                           |                           |+/-1.39E-02    |Jy       |2003AJ....125..525J|1 sigma uncert.        |1.65      microns  |Broad-band measurement                                                                      |061837.71 +782125.3 (J2000)    |Flux integrated from map                                |174.8 x   82.2 arcsec integration area.|From new raw data; Corrected for contaminating sources                                                                                                             
 58    |H (Johnson)         |8.6E+00               |+/-0.03      |mag              |1.82E+14 |4.01E-01    |1.12E-02                  |1.12E-02                  |                           |                           |+/-1.12E-02    |Jy       |1977HarvU.T00M....A|uncertainty            |1.65    microns    |Broad-band measurement                                                                      |                               |Flux in fixed aperture                                  |27.4" aperture                         |From new raw data; derived from a flux in a different bandand a color                                                                                              
 59    |H (Johnson)         |8.2E+00               |+/-0.03      |mag              |1.82E+14 |5.64E-01    |1.58E-02                  |1.58E-02                  |                           |                           |+/-1.58E-02    |Jy       |1977HarvU.T00M....A|uncertainty            |1.65    microns    |Broad-band measurement                                                                      |                               |Flux in fixed aperture                                  |41.1" aperture                         |From new raw data; derived from a flux in a different bandand a color                                                                                              
 60    |H (Johnson)         |7.7E+00               |+/-0.03      |mag              |1.82E+14 |9.28E-01    |2.60E-02                  |2.60E-02                  |                           |                           |+/-2.60E-02    |Jy       |1977HarvU.T00M....A|uncertainty            |1.65    microns    |Broad-band measurement                                                                      |                               |Flux in fixed aperture                                  |105" aperture                          |From new raw data; derived from a flux in a different bandand a color                                                                                              
 61    |K_tot (2MASS LGA)   |7.1E+00               |+/-0.023     |mag              |1.38E+14 |9.97E-01    |2.14E-02                  |2.14E-02                  |                           |                           |+/-2.14E-02    |Jy       |2003AJ....125..525J|1 sigma uncert.        |2.17      microns  |Broad-band measurement                                                                      |061837.71 +782125.3 (J2000)    |Total flux                                              |                                       |From new raw data                                                                                                                                                  
 62    |K_Kron (2MASS LGA)  |7.2E+00               |+/-0.016     |mag              |1.38E+14 |8.90E-01    |1.32E-02                  |1.32E-02                  |                           |                           |+/-1.32E-02    |Jy       |2003AJ....125..525J|1 sigma uncert.        |2.17      microns  |Broad-band measurement                                                                      |061837.71 +782125.3 (J2000)    |Flux integrated from map                                |174.8 x   82.2 arcsec integration area.|From new raw data; Corrected for contaminating sources                                                                                                             
 63    |K_20 (2MASS LGA)    |7.2E+00               |+/-0.016     |mag              |1.38E+14 |9.13E-01    |1.36E-02                  |1.36E-02                  |                           |                           |+/-1.36E-02    |Jy       |2003AJ....125..525J|1 sigma uncert.        |2.17      microns  |Broad-band measurement                                                                      |061837.71 +782125.3 (J2000)    |Flux integrated from map                                |195.0 x   91.7 arcsec integration area.|From new raw data; Corrected for contaminating sources                                                                                                             
 64    |K_s_14arcsec (2MASS)|8.6E+00               |+/-0.015     |mag              |1.38E+14 |2.41E-01    |3.35E-03                  |3.35E-03                  |                           |                           |+/-3.35E-03    |Jy       |20032MASX.C.......:|1 sigma uncert.        |2.17      microns  |Broad-band measurement                                                                      |061837.71 +782125.3 (J2000)    |Flux in fixed aperture                                  |14.0 x 14.0 arcsec aperture            |From new raw data                                                                                                                                                  
 65    |K (Johnson)         |7.7E+00               |+/-0.03      |mag              |1.35E+14 |5.55E-01    |1.55E-02                  |1.55E-02                  |                           |                           |+/-1.55E-02    |Jy       |1977HarvU.T00M....A|uncertainty            |2.22    microns    |Broad-band measurement                                                                      |                               |Flux in fixed aperture                                  |41.1" aperture                         |From new raw data                                                                                                                                                  
 66    |K (Johnson)         |7.2E+00               |+/-0.03      |mag              |1.35E+14 |8.48E-01    |2.37E-02                  |2.37E-02                  |                           |                           |+/-2.37E-02    |Jy       |1977HarvU.T00M....A|uncertainty            |2.22    microns    |Broad-band measurement                                                                      |                               |Flux in fixed aperture                                  |105" aperture                          |From new raw data                                                                                                                                                  
 67    |K (Johnson)         |8.0E+00               |+/-0.03      |mag              |1.35E+14 |4.13E-01    |1.16E-02                  |1.16E-02                  |                           |                           |+/-1.16E-02    |Jy       |1977HarvU.T00M....A|uncertainty            |2.22    microns    |Broad-band measurement                                                                      |                               |Flux in fixed aperture                                  |27.4" aperture                         |From new raw data                                                                                                                                                  
 68    |3.6 microns (IRAC)  |9.5E-01               |+/-2.86E-2   |Jy               |8.44E+13 |9.53E-01    |2.86E-02                  |2.86E-02                  |                           |                           |+/-2.86E-02    |Jy       |2008ApJ...678..804E|rms uncertainty        |3.550 microns      |Broad-band measurement                                                                      |06 18 37.7 +78 21 24.4 (J2000) |Corrected to total flux from single aperture measurement|Color-corrected                        |From new raw data                                                                                                                                                  
 69    |4.5 microns (IRAC)  |7.1E-01               |+/-2.11E-2   |Jy               |6.67E+13 |7.05E-01    |2.11E-02                  |2.11E-02                  |                           |                           |+/-2.11E-02    |Jy       |2008ApJ...678..804E|rms uncertainty        |4.493 microns      |Broad-band measurement                                                                      |06 18 37.7 +78 21 24.4 (J2000) |Corrected to total flux from single aperture measurement|Color-corrected                        |From new raw data                                                                                                                                                  
 71    |5.8 microns (IRAC)  |2.8E+00               |+/-8.49E-2   |Jy               |5.23E+13 |2.83E+00    |8.49E-02                  |8.49E-02                  |                           |                           |+/-8.49E-02    |Jy       |2008ApJ...678..804E|rms uncertainty        |5.731 microns      |Broad-band measurement                                                                      |06 18 37.7 +78 21 24.4 (J2000) |Corrected to total flux from single aperture measurement|Color-corrected                        |From new raw data                                                                                                                                                  
 72    |6 microns (IRS)     |7.4E-01               |             |Jy               |5.00E+13 |7.40E-01    |                          |                          |                           |                           |               |Jy       |2006ApJ...653.1129B|no uncertainty reported|6   microns        |Broad-band measurement                                                                      |06 18 37.71 +78 21 25.3 (J2000)|Flux integrated from map                                |                                       |From new raw data                                                                                                                                                  
 77    |8.0 microns (IRAC)  |9.4E+00               |+/-2.81E-1   |Jy               |3.81E+13 |9.37E+00    |2.81E-01                  |2.81E-01                  |                           |                           |+/-2.81E-01    |Jy       |2008ApJ...678..804E|rms uncertainty        |7.872 microns      |Broad-band measurement                                                                      |06 18 37.7 +78 21 24.4 (J2000) |Corrected to total flux from single aperture measurement|Color-corrected                        |From new raw data                                                                                                                                                  
 82    |12 microns (IRAS)   |7.4E+00               |+/-0.80      |Jy               |2.50E+13 |7.36E+00    |8.00E-01                  |8.00E-01                  |                           |                           |+/-8.00E-01    |Jy       |2004AJ....127.3235S|1 sigma                |12.0   microns     |Broad-band measurement                                                                      |06 10 40.1 +78 22 23 (B1950)   |Flux in fixed aperture                                  |                                       |From reprocessed raw data                                                                                                                                          
 83    |12 microns (IRAS)   |6.8E+00               |+/-0.022     |Jy               |2.50E+13 |6.83E+00    |2.20E-02                  |2.20E-02                  |                           |                           |+/-2.20E-02    |Jy       |2003AJ....126.1607S|1 sigma                |12   microns       |Broad-band measurement                                                                      |06 18 39.8 +78 21 25 (J2000)   |Total flux                                              |Size, Method, Flag codes: MI;see paper |From reprocessed raw data                                                                                                                                          
 84    |12 microns (IRAS)   |6.2E+00               |+/-4   %     |Jy               |2.50E+13 |6.23E+00    |2.49E-01                  |2.49E-01                  |                           |                           |+/-2.49E-01    |Jy       |1990IRASF.C...0000M|uncertainty            |12        microns  |Broad-band measurement                                                                      |061042.3 +782229 (B1950)       |Flux in fixed aperture                                  |IRAS quality flag = 3                  |From new raw data                                                                                                                                                  
 89    |15 microns (IRS)    |2.0E+00               |             |Jy               |2.00E+13 |2.00E+00    |                          |                          |                           |                           |               |Jy       |2006ApJ...653.1129B|no uncertainty reported|15   microns       |Broad-band measurement                                                                      |06 18 37.71 +78 21 25.3 (J2000)|Flux integrated from map                                |                                       |From new raw data                                                                                                                                                  
 94    |24 microns (MIPS)   |1.7E+01               |+/-3.41E-1   |Jy               |1.27E+13 |1.70E+01    |3.41E-01                  |3.41E-01                  |                           |                           |+/-3.41E-01    |Jy       |2008ApJ...678..804E|rms uncertainty        |23.68 microns      |Broad-band measurement                                                                      |06 18 37.7 +78 21 24.4 (J2000) |Corrected to total flux from single aperture measurement|Color-corrected                        |From new raw data                                                                                                                                                  
 95    |25 microns (IRAS)   |2.2E+01               |+/-2.40      |Jy               |1.20E+13 |2.17E+01    |2.40E+00                  |2.40E+00                  |                           |                           |+/-2.40E+00    |Jy       |2004AJ....127.3235S|1 sigma                |25.0   microns     |Broad-band measurement                                                                      |06 10 40.1 +78 22 23 (B1950)   |Flux in fixed aperture                                  |                                       |From reprocessed raw data                                                                                                                                          
 96    |25 microns (IRAS)   |1.9E+01               |+/-0.03      |Jy               |1.20E+13 |1.88E+01    |3.00E-02                  |3.00E-02                  |                           |                           |+/-3.00E-02    |Jy       |2003AJ....126.1607S|1 sigma                |25   microns       |Broad-band measurement                                                                      |06 18 39.8 +78 21 25 (J2000)   |Total flux                                              |Size, Method, Flag codes: MI;see paper |From reprocessed raw data                                                                                                                                          
 97    |25 microns (IRAS)   |1.8E+01               |+/-4   %     |Jy               |1.20E+13 |1.76E+01    |2.49E-01                  |2.49E-01                  |                           |                           |+/-2.49E-01    |Jy       |1990IRASF.C...0000M|uncertainty            |25        microns  |Broad-band measurement                                                                      |061042.3 +782229 (B1950)       |Flux in fixed aperture                                  |IRAS quality flag = 3                  |From new raw data                                                                                                                                                  
 100   |30 microns (IRS)    |2.3E+01               |             |Jy               |9.99E+12 |2.31E+01    |                          |                          |                           |                           |               |Jy       |2006ApJ...653.1129B|no uncertainty reported|30   microns       |Broad-band measurement                                                                      |06 18 37.71 +78 21 25.3 (J2000)|Flux integrated from map                                |                                       |From new raw data                                                                                                                                                  
 104   |52 microns (ISO)    |1.3E+02               |+/-3.2       |Jy               |5.77E+12 |1.35E+02    |3.20E+00                  |3.20E+00                  |                           |                           |+/-3.20E+00    |Jy       |2008ApJS..178..280B|uncertainty            |52 microns         |Broad-band measurement                                                                      |06 18 39.70 +78 21 23.0 (J2000)|Flux integrated from map                                |                                       |From new raw data                                                                                                                                                  
 106   |57 microns (ISO)    |1.6E+02               |+/-2.8       |Jy               |5.26E+12 |1.61E+02    |2.80E+00                  |2.80E+00                  |                           |                           |+/-2.80E+00    |Jy       |2008ApJS..178..280B|uncertainty            |57 microns         |Broad-band measurement                                                                      |06 18 39.70 +78 21 23.0 (J2000)|Flux integrated from map                                |                                       |From new raw data                                                                                                                                                  
 107   |60 microns (IRAS)   |1.5E+02               |+/-16.00     |Jy               |5.00E+12 |1.54E+02    |1.60E+01                  |1.60E+01                  |                           |                           |+/-1.60E+01    |Jy       |2004AJ....127.3235S|1 sigma                |60.0   microns     |Broad-band measurement                                                                      |06 10 40.1 +78 22 23 (B1950)   |Flux in fixed aperture                                  |                                       |From reprocessed raw data                                                                                                                                          
 108   |60 microns (IRAS)   |1.5E+02               |+/-0.063     |Jy               |5.00E+12 |1.47E+02    |6.30E-02                  |6.30E-02                  |                           |                           |+/-6.30E-02    |Jy       |2003AJ....126.1607S|1 sigma                |60   microns       |Broad-band measurement                                                                      |06 18 39.8 +78 21 25 (J2000)   |Total flux                                              |Size, Method, Flag codes: MI;see paper |From reprocessed raw data                                                                                                                                          
 109   |60 microns (ISO)    |1.6E+02               |+/-20  %     |Jy               |5.00E+12 |1.63E+02    |3.27E+01                  |3.27E+01                  |                           |                           |+/-3.27E+01    |Jy       |2001A&A...375..566N|uncertainty            |60   microns       |Broad-band measurement                                                                      |                               |Modelled datum                                          |                                       |From new raw data                                                                                                                                                  
 110   |60 microns (IRAS)   |1.3E+02               |+/-4   %     |Jy               |5.00E+12 |1.31E+02    |5.24E+00                  |5.24E+00                  |                           |                           |+/-5.24E+00    |Jy       |1990IRASF.C...0000M|uncertainty            |60        microns  |Broad-band measurement                                                                      |061042.3 +782229 (B1950)       |Flux in fixed aperture                                  |IRAS quality flag = 3                  |From new raw data                                                                                                                                                  
 111   |63 microns (ISO)    |1.8E+02               |+/-3.2       |Jy               |4.76E+12 |1.83E+02    |3.20E+00                  |3.20E+00                  |                           |                           |+/-3.20E+00    |Jy       |2008ApJS..178..280B|uncertainty            |63 microns         |Broad-band measurement                                                                      |06 18 39.70 +78 21 23.0 (J2000)|Flux integrated from map                                |                                       |From new raw data                                                                                                                                                  
 114   |70 microns (PACS)   |2.0E+02               |+/-0.10E+2   |Jy               |4.28E+12 |1.98E+02    |1.00E+01                  |1.00E+01                  |                           |                           |+/-1.00E+01    |Jy       |2012ApJ...745...95D|uncertainty            |70 microns         |Broad-band measurement                                                                      |06 18 35.6 +78 21 29 (J2000)   |Flux in fixed aperture                                  |                                       |From new raw data                                                                                                                                                  
 115   |70 microns (MIPS)   |1.5E+02               |+/-7.29E+0   |Jy               |4.20E+12 |1.46E+02    |7.29E+00                  |7.29E+00                  |                           |                           |+/-7.29E+00    |Jy       |2008ApJ...678..804E|rms uncertainty        |71.42 microns      |Broad-band measurement                                                                      |06 18 37.7 +78 21 24.4 (J2000) |Corrected to total flux from single aperture measurement|Color-corrected                        |From new raw data                                                                                                                                                  
 116   |88 microns (ISO)    |2.5E+02               |+/-6.2       |Jy               |3.41E+12 |2.50E+02    |6.20E+00                  |6.20E+00                  |                           |                           |+/-6.20E+00    |Jy       |2008ApJS..178..280B|uncertainty            |88 microns         |Broad-band measurement                                                                      |06 18 39.70 +78 21 23.0 (J2000)|Flux integrated from map                                |                                       |From new raw data                                                                                                                                                  
 118   |100 microns (IRAS)  |1.9E+02               |+/-0.24      |Jy               |3.00E+12 |1.94E+02    |2.40E-01                  |2.40E-01                  |                           |                           |+/-2.40E-01    |Jy       |2003AJ....126.1607S|1 sigma                |100   microns      |Broad-band measurement                                                                      |06 18 39.8 +78 21 25 (J2000)   |Total flux                                              |Size, Method, Flag codes: UT;see paper |From reprocessed raw data                                                                                                                                          
 119   |100 microns (IRAS)  |2.2E+02               |+/-24.00     |Jy               |3.00E+12 |2.17E+02    |2.40E+01                  |2.40E+01                  |                           |                           |+/-2.40E+01    |Jy       |2004AJ....127.3235S|1 sigma                |100.0   microns    |Broad-band measurement                                                                      |06 10 40.1 +78 22 23 (B1950)   |Flux in fixed aperture                                  |                                       |From reprocessed raw data                                                                                                                                          
 120   |100 microns (PACS)  |2.3E+02               |+/-0.12E+2   |Jy               |3.00E+12 |2.32E+02    |1.20E+01                  |1.20E+01                  |                           |                           |+/-1.20E+01    |Jy       |2012ApJ...745...95D|uncertainty            |100 microns        |Broad-band measurement                                                                      |06 18 35.6 +78 21 29 (J2000)   |Flux in fixed aperture                                  |                                       |From new raw data                                                                                                                                                  
 121   |100 microns (IRAS)  |1.8E+02               |+/-5   %     |Jy               |3.00E+12 |1.84E+02    |9.21E+00                  |9.21E+00                  |                           |                           |+/-9.21E+00    |Jy       |1990IRASF.C...0000M|uncertainty            |100       microns  |Broad-band measurement                                                                      |061042.3 +782229 (B1950)       |Flux in fixed aperture                                  |IRAS quality flag = 2                  |From new raw data                                                                                                                                                  
 122   |122 microns (ISO)   |1.9E+02               |+/-1.7       |Jy               |2.46E+12 |1.92E+02    |1.70E+00                  |1.70E+00                  |                           |                           |+/-1.70E+00    |Jy       |2008ApJS..178..280B|uncertainty            |122 microns        |Broad-band measurement                                                                      |06 18 39.70 +78 21 23.0 (J2000)|Flux integrated from map                                |                                       |From new raw data                                                                                                                                                  
 124   |145 microns (ISO)   |1.4E+02               |+/-1.8       |Jy               |2.07E+12 |1.39E+02    |1.80E+00                  |1.80E+00                  |                           |                           |+/-1.80E+00    |Jy       |2008ApJS..178..280B|uncertainty            |145 microns        |Broad-band measurement                                                                      |06 18 39.70 +78 21 23.0 (J2000)|Flux integrated from map                                |                                       |From new raw data                                                                                                                                                  
 127   |160 microns (MIPS)  |1.1E+02               |+/-1.35E+1   |Jy               |1.92E+12 |1.12E+02    |1.35E+01                  |1.35E+01                  |                           |                           |+/-1.35E+01    |Jy       |2008ApJ...678..804E|rms uncertainty        |155.90 microns     |Broad-band measurement                                                                      |06 18 37.7 +78 21 24.4 (J2000) |Corrected to total flux from single aperture measurement|Color-corrected                        |From new raw data                                                                                                                                                  
 128   |158 microns (ISO)   |1.4E+02               |+/-4.2       |Jy               |1.90E+12 |1.38E+02    |4.20E+00                  |4.20E+00                  |                           |                           |+/-4.20E+00    |Jy       |2008ApJS..178..280B|uncertainty            |158 microns        |Broad-band measurement                                                                      |06 18 39.70 +78 21 23.0 (J2000)|Flux integrated from map                                |                                       |From new raw data                                                                                                                                                  
 131   |160 microns (PACS)  |1.8E+02               |+/-0.09E+2   |Jy               |1.87E+12 |1.81E+02    |9.00E+00                  |9.00E+00                  |                           |                           |+/-9.00E+00    |Jy       |2012ApJ...745...95D|uncertainty            |160 microns        |Broad-band measurement                                                                      |06 18 35.6 +78 21 29 (J2000)   |Flux in fixed aperture                                  |                                       |From new raw data                                                                                                                                                  
 132   |170 microns (ISO)   |1.2E+02               |+/-3.5       |Jy               |1.76E+12 |1.25E+02    |3.50E+00                  |3.50E+00                  |                           |                           |+/-3.50E+00    |Jy       |2008ApJS..178..280B|uncertainty            |170 microns        |Broad-band measurement                                                                      |06 18 39.70 +78 21 23.0 (J2000)|Flux integrated from map                                |                                       |From new raw data                                                                                                                                                  
 133   |250 microns (SPIRE) |6.6E+01               |+/-0.47E+1   |Jy               |1.20E+12 |6.55E+01    |4.70E+00                  |4.70E+00                  |                           |                           |+/-4.70E+00    |Jy       |2012ApJ...745...95D|uncertainty            |250 microns        |Broad-band measurement                                                                      |06 18 35.6 +78 21 29 (J2000)   |Flux in fixed aperture                                  |                                       |From new raw data                                                                                                                                                  
 134   |350 microns (SPIRE) |2.3E+01               |+/-0.17E+1   |Jy               |8.57E+11 |2.33E+01    |1.70E+00                  |1.70E+00                  |                           |                           |+/-1.70E+00    |Jy       |2012ApJ...745...95D|uncertainty            |350 microns        |Broad-band measurement                                                                      |06 18 35.6 +78 21 29 (J2000)   |Flux in fixed aperture                                  |                                       |From new raw data                                                                                                                                                  
 135   |500 microns (SPIRE) |7.5E+00               |+/-0.53E+0   |Jy               |6.00E+11 |7.45E+00    |5.30E-01                  |5.30E-01                  |                           |                           |+/-5.30E-01    |Jy       |2012ApJ...745...95D|uncertainty            |500 microns        |Broad-band measurement                                                                      |06 18 35.6 +78 21 29 (J2000)   |Flux in fixed aperture                                  |                                       |From new raw data                                                                                                                                                  
 138   |2.8 cm              |3.0E-01               |             |Jy               |1.06E+10 |3.00E-01    |                          |                          |                           |                           |7.00E-02       |Jy       |1973AJ.....78...18M|no uncertainty reported|2.82   cm          |Broad-band measurement                                                                      |061039 +7822 (B1950)           |Integrated from scans                                   |                                       |From new raw data                                                                                                                                                  
 139   |4.5 cm              |3.5E-01               |             |Jy               |6.63E+09 |3.50E-01    |                          |                          |                           |                           |3.00E-02       |Jy       |1973AJ.....78...18M|no uncertainty reported|4.52   cm          |Broad-band measurement                                                                      |061039 +7822 (B1950)           |Integrated from scans                                   |                                       |From new raw data                                                                                                                                                  
 140   |1.49 GHz (VLA)      |1.1E+03               |             |milliJy          |1.49E+09 |1.07E+00    |                          |                          |                           |                           |               |Jy       |1996ApJS..103...81C|no uncertainty reported|1.49   GHz         |Broad-band measurement                                                                      |061040.3 +782228 (B1950)       |Flux integrated from map                                |Beamwidth = 60"                        |Averaged from previously published data                                                                                                                            
 141   |1.49 GHz (VLA)      |1.1E+03               |             |milliJy          |1.49E+09 |1.09E+00    |                          |                          |                           |                           |               |Jy       |1996ApJS..103...81C|no uncertainty reported|1.490   GHz        |Broad-band measurement                                                                      |061040.8 +782227 (B1950)       |Total flux                                              |Beamwidth = 60"                        |Averaged from previously published data                                                                                                                            
 142   |1465 MHz            |1.0E+03               |+/-40        |milliJy          |1.46E+09 |1.02E+00    |4.00E-02                  |4.00E-02                  |                           |                           |+/-4.00E-02    |Jy       |1983ApJS...53..459C|rms uncertainty        |1465       MHz     |Broad-band measurement                                                                      |                               |Flux integrated from map                                |                                       |From new raw data                                                                                                                                                  
 148   |1.4GHz              |1.1E+03               |+/-40.0      |milliJy          |1.40E+09 |1.07E+00    |4.00E-02                  |4.00E-02                  |                           |                           |+/-4.00E-02    |Jy       |1998AJ....115.1693C|uncertainty            |1.40   GHz         |Broad-band measurement                                                                      |06 18 37.71 +78 21 23.9 (J2000)|Flux integrated from map                                |                                       |From new raw data                                                                                                                                                  
 149   |1.40 GHz            |1.2E+03               |             |milliJy          |1.40E+09 |1.23E+00    |                          |                          |                           |                           |               |Jy       |1992ApJS...79..331W|no uncertainty reported|1.4        GHz     |Broad-band measurement                                                                      |061033.6 +782120 (B1950)       |Flux integrated from map                                |                                       |From new raw data                                                                                                                                                  
 150   |1400 MHz (NRAO)     |1.3E+00               |             |Jy               |1.40E+09 |1.30E+00    |                          |                          |                           |                           |               |Jy       |1964AJ.....69..277H|no uncertainty reported|1400      MHz      |Broad-band measurement; peak value reported                                                 |061039 +7824 (B1950)           |Peak flux                                               |                                       |From new raw data                                                                                                                                                  
 151   |1.4 GHz (VLA)       |1.1E+03               |             |milliJy          |1.40E+09 |1.07E+00    |                          |                          |                           |                           |               |Jy       |2002AJ....124..675C|no uncertainty reported|1.4   GHz          |Broad-band measurement                                                                      |                               |Flux integrated from map                                |                                       |Averaged from previously published data                                                                                                                            
 152   |1365 MHz (WSRT)     |1.1E+03               |+/-10        |milliJy          |1.37E+09 |1.10E+00    |1.00E-02                  |1.00E-02                  |                           |                           |+/-1.00E-02    |Jy       |2007A&A...461..455B|uncertainty            |1365   MHz         |Broad-band measurement                                                                      |                               |Total flux                                              |                                       |From new raw data                                                                                                                                                  
 153   |750 MHz (NRAO)      |1.6E+00               |             |Jy               |7.50E+08 |1.60E+00    |                          |                          |                           |                           |               |Jy       |1964AJ.....69..277H|no uncertainty reported|750      MHz       |Broad-band measurement; peak value reported                                                 |061039 +7824 (B1950)           |Peak flux                                               |                                       |From new raw data                                                                                                                                                  
 154   |92 cm (WENSS)       |2.0E+03               |+/-82.0      |milliJy          |3.52E+08 |2.05E+00    |8.20E-02                  |8.20E-02                  |                           |                           |+/-8.20E-02    |Jy       |1998WENSP.C.......:|uncertainty            |92         cm      |Broad-band measurement                                                                      |061039.79 +782227.7 (B1950)    |Peak flux                                               |Single component source                |From new raw data                                                                                                                                                  
 155   |92 cm (WENSS)       |2.5E+03               |+/-100.5     |milliJy          |3.52E+08 |2.51E+00    |1.00E-01                  |1.00E-01                  |                           |                           |+/-1.00E-01    |Jy       |1998WENSP.C.......:|uncertainty            |92         cm      |Broad-band measurement                                                                      |061039.79 +782227.7 (B1950)    |Flux integrated from map                                |Single component source                |From new raw data                                                                                                                                                  
 156   |178 MHz             |3.2E+00               |+/-15.0%     |Jy               |1.78E+08 |3.20E+00    |4.80E-01                  |4.80E-01                  |                           |                           |+/-4.80E-01    |Jy       |1967MmRAS..71...49G|uncertainty            |178        MHz     |Broad-band measurement                                                                      |061040.1 +782012 (B1950)       |Integrated from scans                                   |                                       |From new raw data; Uncorrected for known sources in beam                                                                                                           
 157   |151 MHz (6C)        |4.0E+00               |+/-0.090     |Jy               |1.52E+08 |4.04E+00    |9.00E-02                  |9.00E-02                  |                           |                           |+/-9.00E-02    |Jy       |1991MNRAS.251...46H|typical accuracy       |151.5      MHz     |Broad-band measurement                                                                      |061040.6 782232. (B1950)       |Flux integrated from map                                |                                       |From new raw data                                                                                                                                                  
 158   |151 MHz (6C)        |3.7E+00               |+/-0.040     |Jy               |1.52E+08 |3.73E+00    |4.00E-02                  |4.00E-02                  |                           |                           |+/-4.00E-02    |Jy       |1991MNRAS.251...46H|typical accuracy       |151.5      MHz     |Broad-band measurement                                                                      |061040.6 782232. (B1950)       |Peak flux                                               |                                       |From new raw data                                                                                                                                                  
 159   |74 MHz (VLA)        |4.2E+00               |+/-0.45      |Jy               |7.38E+07 |4.21E+00    |4.50E-01                  |4.50E-01                  |                           |                           |+/-4.50E-01    |Jy       |2007AJ....134.1245C|rms uncertainty        |73.8   MHz         |Broad-band measurement                                                                      |06 18 37.55 +78 21 21.7 (J2000)|Flux integrated from map                                |Corrected for clean bias               |From new raw data                                                                                                                                                  
 160   |57.5 MHz            |6.9E+00               |+/-1.7       |Jy               |5.75E+07 |6.90E+00    |1.70E+00                  |1.70E+00                  |                           |                           |+/-1.70E+00    |Jy       |1990ApJ...352...30I|uncertainty            |57.5       MHz     |Broad-band measurement                                                                      |                               |Flux integrated from map                                |                                       |From new raw data                                                                                                                                                  
 161   |38 MHz (8C)         |8.1E+00               |+/-0.8       |Jy               |3.78E+07 |8.10E+00    |8.33E-01                  |8.33E-01                  |                           |                           |+/-8.33E-01    |Jy       |1995MNRAS.274..447H|2.5 times noise        |38         MHz     |Broad-band measurement                                                                      |061036. +782233. (B1950)       |Flux integrated from map                                |Single component source                |From new raw data                                                                                                                                                  
 162   |38 MHz (8C)         |5.8E+00               |+/-15.0%     |Jy               |3.78E+07 |5.80E+00    |8.70E-01                  |8.70E-01                  |                           |                           |+/-8.70E-01    |Jy       |1995MNRAS.274..447H|no uncertainty reported|38         MHz     |Broad-band measurement                                                                      |061036. +782233. (B1950)       |Peak flux                                               |Single component source                |From new raw data                                                                                                                                                  
