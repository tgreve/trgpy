
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-04-05T08:15:36PDT



Photometric Data for SDSS J163655.77+405910.0

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|2-8 keV (Chandra)   | 1.47E-14  |+/-0.21E-14|ergs cm^-2^ s^-1^   |1.21E+18|  1.22E-09|+/-1.74E-10|Jy|2003MNRAS.343..293M|uncertainty|       5   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
2|0.5-8 keV (Chandra) | 1.02E-14  |+/-0.11E-14|ergs cm^-2^ s^-1^   |1.03E+18|  9.93E-10|+/-1.07E-10|Jy|2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
3|0.5-2 keV (Chandra) | 0.21E-14  |+/-0.04E-14|ergs cm^-2^ s^-1^   |3.02E+17|  6.95E-10|+/-1.32E-10|Jy|2003MNRAS.343..293M|uncertainty|    1.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
4|U_aper_ (INT/WFC)   | 22.63     |+/-0.10 |mag                 |8.37E+14|  1.37E-06|+/-1.26E-07|Jy|2005MNRAS.358..333G|uncertainty|    3581   A         | Broad-band measurement|249.23262 +40.98589 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data
5|[O II] 3727 (SUBARU)| 3.6E-16   |+/-0.9E-16|ergs cm^-2^ s^-1^   |8.04E+14|  4.48E-08|+/-1.12E-08|Jy|2006ApJ...651..713T|uncertainty|    3727   A         | Line measurement; flux integrated over line; lines measured in emission| | Flux integrated from map|                                        |From new raw data
6|g'_aper_ (INT/WFC)  | 22.87     |+/-0.04 |mag                 |6.19E+14|  2.79E-06|+/-1.03E-07|Jy|2005MNRAS.358..333G|uncertainty|    4846   A         | Broad-band measurement|249.23262 +40.98589 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data
7|H{beta} (SUBARU)    | 2.7E-16   |+/-1.0E-16|ergs cm^-2^ s^-1^   |6.17E+14|  4.38E-08|+/-1.62E-08|Jy|2006ApJ...651..713T|uncertainty|    4861   A         | Line measurement; flux integrated over line; lines measured in emission| | Flux integrated from map|                                        |From new raw data
8|[O III] 4959 SUBARU | 15.7E-16  |+/-1.6E-16|ergs cm^-2^ s^-1^   |6.05E+14|  2.60E-07|+/-2.64E-08|Jy|2006ApJ...651..713T|uncertainty|    4959   A         | Line measurement; flux integrated over line; lines measured in emission| | Flux integrated from map|                                        |From new raw data
9|[O III] 5007 SUBARU | 47.1E-16  |+/-1.6E-16|ergs cm^-2^ s^-1^   |5.99E+14|  7.86E-07|+/-2.67E-08|Jy|2006ApJ...651..713T|uncertainty|    5007   A         | Line measurement; flux integrated over line; lines measured in emission| | Flux integrated from map|                                        |From new raw data
10|r'_tot_ (INT/WFC)   | 23.09     |+/-0.11 |mag                 |4.80E+14|  1.81E-06|+/-1.84E-07|Jy|2005MNRAS.358..333G|uncertainty|    6240   A         | Broad-band measurement|249.23262 +40.98589 (J2000)| Total flux|                                        |Averaged new and previously published data
11|r'_aper_ (INT/WFC)  | 22.92     |+/-0.08 |mag                 |4.80E+14|  2.12E-06|+/-1.56E-07|Jy|2005MNRAS.358..333G|uncertainty|    6240   A         | Broad-band measurement|249.23262 +40.98589 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data
12|H{alpha} (SUBARU)   | 18.4E-16  |+/-2.4E-16|ergs cm^-2^ s^-1^   |4.57E+14|  4.03E-07|+/-5.25E-08|Jy|2006ApJ...651..713T|uncertainty|    6563   A         | Line measurement; flux integrated over line; lines measured in emission| | Flux integrated from map|                                        |From new raw data
13|H{alpha} (Keck)     | 2.4E-19   |+/-0.4E-19| W/m^2^             |4.57E+14|  5.25E-08|+/-8.75E-09|Jy|2004ApJ...617...64S|uncertainty|      6563 A         | Line measurement; flux integrated over line; lines measured in emission|163655.80 +405914.0 (J2000)| Flux integrated from map|                                        |From new raw data
14|H{alpha} (Keck)     | 16E-19    |+/-2E-19| W/m^2^             |4.57E+14|  3.50E-07|+/-4.38E-08|Jy|2004ApJ...617...64S|uncertainty|      6563 A         | Line measurement; flux integrated over line; lines measured in emission|163655.80 +405914.0 (J2000)| Flux integrated from map|Broad-line component                    |From new raw data
15|i'_aper_ (INT/WFC)  | 23.02     |+/-0.23 |mag                 |3.87E+14|  1.56E-06|+/-3.29E-07|Jy|2005MNRAS.358..333G|uncertainty|    7743   A         | Broad-band measurement|249.23262 +40.98589 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data
16|I (Cousins)         | |>25.90     |mag                 |3.79E+14| |1.11E-07|Jy|2004ApJ...616...71S|3sigma uncertainty|    7900   A         | Broad-band measurement| | Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
17|K_s_ (2MASS)        | |>20.50     |mag                 |1.38E+14| |4.21E-06|Jy|2004ApJ...616...71S|3sigma uncertainty|    2.17   microns   | Broad-band measurement| | Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
18|2.2 microns (IRS)   | 0.387     |+/-0.009| milliJy            |1.36E+14|  3.87E-04|+/-9.00E-06|Jy|2009MNRAS.395.1695H|uncertainty|       2.2 microns   | Broad-band measurement| | Flux in fixed aperture|                                        |From new raw data
19|3.6 microns (IRAC)  | 27.580    |+/-0.520| microJy            |8.44E+13|  2.76E-05|+/-5.20E-07|Jy|2009AJ....137.3884R|uncertainty|     3.550 microns   | Broad-band measurement|249.232388 40.986118 (J2000)| Flux integrated from map|                                        |From new raw data
20|3.6 microns (IRAC)  | 27.6      |+/-0.5  | microJy            |8.44E+13|  2.76E-05|+/-5.00E-07|Jy|2009MNRAS.395.1695H|uncertainty|     3.550 microns   | Broad-band measurement| | Flux in fixed aperture|                                        |From new raw data
21|4.5 microns (IRAC)  | 52.640    |+/-0.960| microJy            |6.67E+13|  5.26E-05|+/-9.60E-07|Jy|2009AJ....137.3884R|uncertainty|     4.493 microns   | Broad-band measurement|249.232388 40.986118 (J2000)| Flux integrated from map|                                        |From new raw data
22|4.5 microns (IRAC)  | 52.6      |+/-1.0  | microJy            |6.67E+13|  5.26E-05|+/-1.00E-06|Jy|2009MNRAS.395.1695H|uncertainty|     4.493 microns   | Broad-band measurement| | Flux in fixed aperture|                                        |From new raw data
23|5.5 microns (IRS)   | 2.33      |+/-0.25 | milliJy            |5.45E+13|  2.33E-03|+/-2.50E-04|Jy|2009MNRAS.395.1695H|uncertainty|       5.5 microns   | Broad-band measurement| | Flux in fixed aperture|                                        |From new raw data
24|5.8 microns (IRAC)  | 120.700   |+/-3.590| microJy            |5.23E+13|  1.21E-04|+/-3.59E-06|Jy|2009AJ....137.3884R|uncertainty|     5.731 microns   | Broad-band measurement|249.232388 40.986118 (J2000)| Flux integrated from map|                                        |From new raw data
25|5.8 microns (IRAC)  | 121       |+/-3    | microJy            |5.23E+13|  1.21E-04|+/-3.00E-06|Jy|2009MNRAS.395.1695H|uncertainty|     5.731 microns   | Broad-band measurement| | Flux in fixed aperture|                                        |From new raw data
26|7 microns (IRS)     | 2.7       |+/-0.2  | milliJy            |4.28E+13|  2.70E-03|+/-2.00E-04|Jy|2009MNRAS.395.1695H|uncertainty|         7 microns   | Broad-band measurement| | Flux in fixed aperture|                                        |From new raw data
27|8.0 microns (IRAC)  | 398.910   |+/-4.250| microJy            |3.81E+13|  3.99E-04|+/-4.25E-06|Jy|2009AJ....137.3884R|uncertainty|     7.872 microns   | Broad-band measurement|249.232388 40.986118 (J2000)| Flux integrated from map|                                        |From new raw data
28|8.0 microns (IRAC)  | 399       |+/-4    | microJy            |3.81E+13|  3.99E-04|+/-4.00E-06|Jy|2009MNRAS.395.1695H|uncertainty|     7.872 microns   | Broad-band measurement| | Flux in fixed aperture|                                        |From new raw data
30|15 microns (IRS)    | 8.3       |+/-1.3  | milliJy            |2.00E+13|  8.30E-03|+/-1.30E-03|Jy|2009MNRAS.395.1695H|uncertainty|        15 microns   | Broad-band measurement| | Flux in fixed aperture|                                        |From new raw data
31|24 microns (MIPS)   | 2.39      |+/-0.02 | milliJy            |1.27E+13|  2.39E-03|+/-2.00E-05|Jy|2009MNRAS.395.1695H|uncertainty|     23.68 microns   | Broad-band measurement| | Flux in fixed aperture|                                        |From new raw data
32|70 microns (MIPS)   | 13.0      |+/-1.2  | milliJy            |4.20E+12|  1.30E-02|+/-1.20E-03|Jy|2009MNRAS.395.1695H|uncertainty|     71.42 microns   | Broad-band measurement| | Flux in fixed aperture|                                        |From new raw data
33|850 microns (SCUBA) | -0.5      |+/-1.4  | milliJy            |3.53E+11|-0.5E-03 |+/-1.40E-03|Jy|2004ApJ...614..671C|1 sigma|       850 microns   | Broad-band measurement|163656.28 +405912.2 (J2000)| Flux integrated from map|                                        |From new raw data
34|850 microns (SCUBA) | 8.7       |+/-2.1  | milliJy            |3.53E+11|8.7E-03|+/-2.1E-03|Jy|2004ApJ...614..671C|1 sigma|       850 microns   | Broad-band measurement|163656.28 +405912.2 (J2000)| Flux integrated from map|                                        |From new raw data
35|1200 microns (MAMBO)| 2.2       |+/-0.6  | milliJy            |2.50E+11|  2.20E-03|+/-6.00E-04|Jy|2004MNRAS.354..779G|uncertainty|      1200 microns   | Broad-band measurement|16 36 55.9 +40 59 12 (J2000)| Flux integrated from map|S/N = 3.66                              |From new raw data
36|1.4 GHz (VLA)       | 200       |+/-23   | microJy            |1.40E+09|  2.00E-04|+/-2.30E-05|Jy|2006MNRAS.371..963B|1 sigma|       1.4 GHz       | Broad-band measurement|16 36 55.767 +40 59 09.97 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
