
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-05-28T01:42:09PDT



Photometric Data for LABd05, z=2.656

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|3.6 microns (IRAC)  | 20.4      |+/-2.6  |microJy             |8.44E+13|  2.04E-05|+/-2.60E-06|Jy|2012ApJ...744..150B|uncertainty|     3.550 microns   | Broad-band measurement|218.545783 +33.292419 (J2000)| Corrected to total flux from single aperture measurement|                                        |From reprocessed raw data
2|4.5 microns (IRAC)  | 26.3      |+/-3.1  |microJy             |6.67E+13|  2.63E-05|+/-3.10E-06|Jy|2011ApJ...728...59C|uncertainty|     4.493 microns   | Broad-band measurement|| Flux in fixed aperture|                                        |From reprocessed raw data
3|4.5 microns (IRAC)  | 26.3      |+/-3.4  |microJy             |6.67E+13|  2.63E-05|+/-3.40E-06|Jy|2012ApJ...744..150B|uncertainty|     4.493 microns   | Broad-band measurement|218.545783 +33.292419 (J2000)| Corrected to total flux from single aperture measurement|                                        |From reprocessed raw data
4|5.8 microns (IRAC)  | 49.7      |+/-16.9 |microJy             |5.23E+13|  4.97E-05|+/-1.69E-05|Jy|2012ApJ...744..150B|uncertainty|     5.731 microns   | Broad-band measurement|218.545783 +33.292419 (J2000)| Corrected to total flux from single aperture measurement|                                        |From reprocessed raw data
5|8.0 microns (IRAC)  | 77.0      |+/-14.9 |microJy             |3.81E+13|  7.70E-05|+/-1.49E-05|Jy|2011ApJ...728...59C|uncertainty|     7.872 microns   | Broad-band measurement|| Flux in fixed aperture|                                        |From reprocessed raw data
6|8.0 microns (IRAC)  | 76.9      |+/-15.0 |microJy             |3.81E+13|  7.69E-05|+/-1.50E-05|Jy|2012ApJ...744..150B|uncertainty|     7.872 microns   | Broad-band measurement|218.545783 +33.292419 (J2000)| Corrected to total flux from single aperture measurement|                                        |From reprocessed raw data
7|24 microns (MIPS)   | 860       |+/-50   |microJy             |1.27E+13|  8.60E-04|+/-5.00E-05|Jy|2011ApJ...728...59C|uncertainty|     23.68 microns   | Broad-band measurement|| Flux integrated from map|                                        |From reprocessed raw data
8|24 microns (MIPS)   | 860       |+/-51   |microJy             |1.27E+13|  8.60E-04|+/-5.10E-05|Jy|2012ApJ...744..150B|uncertainty|     23.68 microns   | Broad-band measurement|218.545783 +33.292419 (J2000)| Corrected to total flux from single aperture measurement|                                        |From reprocessed raw data
9|70 microns (MIPS)   ||<9         |milliJy             |4.20E+12||9.00E-03|Jy|2012ApJ...744..178Y|3 sigma|     71.42 microns   | Broad-band measurement|14 34 11.0 33 17 33 (J2000)| Flux in fixed aperture|                                        |From new raw data
10|160 microns (MIPS)  ||<51        |milliJy             |1.92E+12||5.10E-02|Jy|2012ApJ...744..178Y|3 sigma|     155.9 microns   | Broad-band measurement|14 34 11.0 33 17 33 (J2000)| Flux in fixed aperture|                                        |From new raw data
11|250 microns (SPIRE  | 18.8      |+/-5.2  |milliJy             |1.20E+12|  1.88E-02|+/-5.20E-03|Jy|2012ApJ...744..178Y|uncertainty|       250 microns   | Broad-band measurement|14 34 11.0 33 17 33 (J2000)| Flux in fixed aperture|                                        |From new raw data
12|350 microns SHARC-II| 37        |+/-13   |milliJy             |8.57E+11|  3.70E-02|+/-1.30E-02|Jy|2009ApJ...705..184B|uncertainty|       350 microns   | Broad-band measurement|14 34 10.980 +33 17 32.70 (J2000)| Flux in fixed aperture|20" diameter aperture                   |From new raw data
13|350 microns (SPIRE  | 26.9      |+/-5.1  |milliJy             |8.57E+11|  2.69E-02|+/-5.10E-03|Jy|2012ApJ...744..178Y|uncertainty|       350 microns   | Broad-band measurement|14 34 11.0 33 17 33 (J2000)| Flux in fixed aperture|                                        |From new raw data
14|1200 microns (MAMBO) | 2.76      |+/-0.35 |milliJy             |2.50E+11|  2.76E-03|+/-3.50E-04|Jy|2012ApJ...744..178Y|uncertainty|      1200 microns   | Broad-band measurement|14 34 11.0 33 17 33 (J2000)| Flux in fixed aperture|                                        |From new raw data
1|1900 microns (PdBI)   | 0.38   | 0.05   |mJy                 |1.576215e+11 |0.38E-03 |+/-0.05E-03|Jy|2010ApJ...709..210K|3sigma uncertainty|      1900  microns   | Broad-band measurement|16 35 55.67 +66 12 59.51 (J2000)| Flux integrated from map|                                        |From new raw data
2|3169 microns (PdBI)   ||<0.15   |mJy                 |9.45831E+10|         |0.15E-03|Jy|2010ApJ...709..210K|3sigma uncertainty|      3169  microns   | Broad-band measurement|16 35 55.67 +66 12 59.51 (J2000)| Flux integrated from map|                                        |From new raw data
15|1.38 GHz (WSRT)     | 0.14      |+/-0.04 | milliJy            |1.38E+09|  1.40E-04|+/-4.00E-05|Jy|2002AJ....123.1784D|uncertainty|      1.38 GHz       | Broad-band measurement|218.5449 +33.2909 (J2000)| Flux integrated from map|a = 0"; b = 0"; PA = 0 deg              |From new raw data
