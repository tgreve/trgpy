\queryDateTime = 2019-01-31T03:55:18PST
\Description = Published and Homogenized [Frequency, Flux Dens...
\source = /local/home/nedops/pkgs/apache-tomcat-7.0.82/temp/workarea/firefly/temp_files/IpacTableFromSource1734216149608410155.tbl
\LINK = http://ned.ipac.caltech.edu/cgi-bin/datasearch?sea
\QUERY_STATUS = OK
\CatalogTargetColName = Coordinates Targeted
\tblFilePath = ${temp-files}/89A/IpacTableFromSource_ddac4e29eeefa15fc4be86febae672a8.hsql
\title = photandseds
\resultSetID = data_a2fda9d5438748ff3127079c32ca8ff0
\resultSetRequest = {"RequestClass":"ServerRequest","META_INFO":{"tblFilePath":"${temp-files}\/FDE\/IpacTableFromSource_f5895644fd2b25addc26423e2cebd560.hsql","col.Upper limit of uncertainty.PrefWidth":"10","col.Spatial Mode.PrefWidth":"22","col.Refcode.FmtDisp":"<a HREF=\"javascript:getReferenceInfo('%s','_nedInternal');\">&nbsp;&nbsp;&nbsp;Ref &swarr;<\/a>","col.Units.PrefWidth":"6","col.Flux Density.FmtDisp":"%e","title":"photandseds","col.Qualifiers.PrefWidth":"22","col.Significance.PrefWidth":"16","col.Coordinates Targeted.PrefWidth":"24","tblFileType":"hsql","tbl_id":"tbl_id-c7911-19","col.Lower limit of uncertainty.PrefWidth":"10","col.Photometry Measurement.FmtDisp":"%e","col.Lower limit of Flux Density.PrefWidth":"10","col.Frequency Mode.PrefWidth":"22","col.Comments.PrefWidth":"26","col.Upper limit of Flux Density.PrefWidth":"10","col.Refcode.PrefWidth":"8"},"tbl_id":"tbl_id-c7911-19","startIdx":0,"pageSize":500,"alt_source":"http:\/\/ned.ipac.caltech.edu\/cgi-bin\/datasearch?meas_type=bot&ebars_spec=ebars&label_spec=no&x_spec=freq&y_spec=Fnu_jy&xr=-1&of=xml_main&search_type=Photometry&objname=ngc1365&hconst=67.8&omegam=0.308&omegav=0.692&corr_z=1","id":"IpacTableFromSource","source":"http:\/\/ned.ipac.caltech.edu\/cgi-bin\/datasearch?meas_type=bot&ebars_spec=ebars&label_spec=no&x_spec=freq&y_spec=Fnu_jy&xr=-1&of=xml_main&search_type=Photometry&objname=ngc1365&hconst=67.8&omegam=0.308&omegav=0.692&corr_z=1","filters":"\"NED Units\" = 'Jy'"}
\tblFileType = hsql
\tbl_id = tbl_id-c7911-19
\
z=0.00546
|No.|Observed Passband   |Photometry Measurement|Uncertainty |Units               |Frequency|Flux Density|Upper limit of uncertainty|Lower limit of uncertainty|Upper limit of Flux Density|Lower limit of Flux Density|NED Uncertainty|NED Units|Refcode                                                                                                       |Significance           |Published frequency|Frequency Mode                                                         |Coordinates Targeted             |Spatial Mode                                             |Qualifiers                              |Comments                                                                                                                                                           |
|int|char                |double                |char        |char                |double   |double      |double                    |double                    |double                     |double                     |char           |char     |char                                                                                                          |char                   |char               |char                                                                   |char                             |char                                                     |char                                    |char                                                                                                                                                               |
|   |                    |                      |            |                    |Hz       |Jy          |                          |                          |                           |                           |               |         |                                                                                                              |                       |                   |                                                                       |                                 |                                                         |                                        |                                                                                                                                                                   |
|   |                    |                      |            |                    |         |            |                          |                          |                           |                           |               |         |                                                                                                              |                       |                   |                                                                       |                                 |                                                         |                                        |                                                                                                                                                                   |
   1|14-195 keV (Swift)  |          7.190000e-11|+/-0.44E-11 |erg/s/cm^2^         | 2.53E+19|2.840000e-07|                  1.74E-08|                  1.74E-08|                           |                           |+/-1.74E-08    |Jy       |<a HREF="javascript:getReferenceInfo('2010ApJS..186..378T','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |104.50 keV         |Broad-band measurement                                                 |053.377 -36.111 (J2000)          |Flux integrated from map                                 |                                        |From new raw data; NED frequency assigned to mid-point ofband in keV                                                                                               
   2|14-195 keV (Swift)  |          7.200000e-11|            |erg/cm^2^/s         | 2.53E+19|2.850000e-07|                          |                          |                           |                           |               |Jy       |<a HREF="javascript:getReferenceInfo('2008ApJ...681..113T','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|104.50 keV         |Broad-band measurement                                                 |053.4015 -36.1404 (J2000)        |Modelled datum                                           |                                        |From new raw data; NED frequency assigned to mid-point ofband in keV                                                                                               
   3|15-150 keV (Swift)  |          5.600000e-11|+/-3.2e-12  |erg/cm^2^/s         | 1.99E+19|2.810000e-07|                  1.61E-08|                  1.61E-08|                           |                           |+/-1.61E-08    |Jy       |<a HREF="javascript:getReferenceInfo('2010A&A...524A..64C','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |82.50 keV          |Broad-band measurement                                                 |053.381 -36.143 (J2000)          |Modelled datum                                           |                                        |From new raw data; NED frequency assigned to mid-point ofband in keV                                                                                               
   4|40-100 keV INTEGRAL |          2.200000e-11|            |erg/cm^2^/s         | 1.69E+19|1.300000e-07|                          |                          |                           |                           |               |Jy       |<a HREF="javascript:getReferenceInfo('2009A&A...505..417B','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|70.00 keV          |Broad-band measurement                                                 |53.40208 -36.13806 (J2000)       |Modelled datum                                           |                                        |From new raw data; NED frequency assigned to mid-point ofband in keV                                                                                               
   5|20-100 keV (Suzaku) |          7.200000e-11|            |erg/s/cm^2^         | 1.45E+19|4.970000e-07|                          |                          |                           |                           |               |Jy       |<a HREF="javascript:getReferenceInfo('2009ApJ...705L...1R','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|60.00 keV          |Broad-band measurement                                                 |                                 |Modelled datum                                           |Observed flux                           |From new raw data; NED frequency assigned to mid-point ofband in keV                                                                                               
   6|17-60 keV (INTEGRAL)|          3.300000e-11|+/-0.65E-11 |erg s^-1^ cm^-2^    | 9.31E+18|3.540000e-07|                  6.98E-08|                  6.98E-08|                           |                           |+/-6.98E-08    |Jy       |<a HREF="javascript:getReferenceInfo('2007A&A...462...57S','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |38.50   keV        |Broad-band measurement                                                 |                                 |Flux integrated from map                                 |                                        |Averaged new and previously published data; NED frequencyassigned to mid-point of band in keV                                                                      
   7|15-55 keV (Swift)   |          3.120000e-11|+/-0.17E-11 |erg/cm^2^/s         | 8.46E+18|3.690000e-07|                  2.01E-08|                  2.01E-08|                           |                           |+/-2.01E-08    |Jy       |<a HREF="javascript:getReferenceInfo('2009ApJ...699..603A','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |35.00 keV          |Broad-band measurement                                                 |053.433 -36.141 (J2000)          |Flux integrated from map                                 |                                        |From reprocessed raw data; NED frequency assigned tomid-point of band in keV                                                                                       
   8|20-40 keV (INTEGRAL)|          1.500000e-11|            |erg/cm^2^/s         | 7.25E+18|2.070000e-07|                          |                          |                           |                           |               |Jy       |<a HREF="javascript:getReferenceInfo('2009A&A...505..417B','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|30.00 keV          |Broad-band measurement                                                 |53.40208 -36.13806 (J2000)       |Modelled datum                                           |                                        |From new raw data; NED frequency assigned to mid-point ofband in keV                                                                                               
   9|20-40 keV (INTEGRAL)|          2.100000e-11|+/-0.876E-11|erg/s/cm^2^         | 7.25E+18|2.900000e-07|                  1.21E-07|                  1.21E-07|                           |                           |+/-1.21E-07    |Jy       |<a HREF="javascript:getReferenceInfo('2010A&A...522A..68T','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|2 sigma                |30.00 keV          |Broad-band measurement                                                 |                                 |Flux integrated from map                                 |                                        |From new raw data; NED frequency assigned to mid-point ofband in keV                                                                                               
  10|10-50 keV (Suzaku)  |          1.770000e+00|            |log(erg/s/cm^2^)    | 7.25E+18|8.120000e-07|                          |                          |                           |                           |               |Jy       |<a HREF="javascript:getReferenceInfo('2011ApJ...727...19F','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|30.00 keV          |Broad-band measurement                                                 |                                 |Modelled datum                                           |                                        |From reprocessed raw data; NED frequency assigned tomid-point of band in keV                                                                                       
  11|2-10 keV            |          6.600000e-15|            |W/m^2^              | 1.45E+18|4.550000e-07|                          |                          |                           |                           |4.55E-07       |Jy       |<a HREF="javascript:getReferenceInfo('2004A&A...418..465L','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|6   keV            |Broad-band measurement                                                 |                                 |Flux integrated from map                                 |Observed flux                           |Averaged from previously published data; NED frequencyassigned to mid-point of band in keV                                                                         
  12|2-10 keV            |          2.310000e-14|            |W/m^2^              | 1.45E+18|1.590000e-06|                          |                          |                           |                           |               |Jy       |<a HREF="javascript:getReferenceInfo('2004A&A...418..465L','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|6   keV            |Broad-band measurement                                                 |                                 |Flux integrated from map                                 |Intrinsic flux                          |Averaged from previously published data; Extinction-correctedfor Milky Way; NED frequency assigned to mid-point of band in keV                                     
  13|2-10 keV (Swift)    |          8.800000e-13|            |erg/s/cm^2^         | 1.45E+18|6.070000e-08|                          |                          |                           |                           |               |Jy       |<a HREF="javascript:getReferenceInfo('2009ApJ...690.1322W','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|6.00 keV           |Broad-band measurement                                                 |03 33 36.4 -36 08 25.4 (J2000)   |Modelled datum                                           |                                        |From new raw data; NED frequency assigned to mid-point ofband in keV                                                                                               
  14|2-10 keV (XMM)      |          1.370000e-11|            |erg/s/cm^2^         | 1.45E+18|9.450000e-07|                          |                          |                           |                           |               |Jy       |<a HREF="javascript:getReferenceInfo('2009ApJ...696..160R','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|6.00 keV           |Broad-band measurement                                                 |                                 |Flux integrated from map                                 |Observed flux                           |From new raw data; NED frequency assigned to mid-point ofband in keV                                                                                               
  15|2-10 keV (Suzaku)   |          1.300000e-11|            |erg/s/cm^2^         | 1.45E+18|8.970000e-07|                          |                          |                           |                           |               |Jy       |<a HREF="javascript:getReferenceInfo('2009ApJ...705L...1R','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|6.00 keV           |Broad-band measurement                                                 |                                 |Modelled datum                                           |Observed flux                           |From new raw data; NED frequency assigned to mid-point ofband in keV                                                                                               
  16|2-10 keV (XMM)      |          1.300000e-11|            |erg/s/cm^2^         | 1.45E+18|8.940000e-07|                          |                          |                           |                           |               |Jy       |<a HREF="javascript:getReferenceInfo('2011MNRAS.413.1206B','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|6.00 keV           |Broad-band measurement                                                 |053.402 -36.140 (J2000)          |Modelled datum                                           |                                        |From reprocessed raw data; NED frequency assigned tomid-point of band in keV                                                                                       
  17|0.5-10 keV (Suzaku) |          1.280000e-11|+/-0.83E-12 |erg/cm^2^/s         | 1.27E+18|1.010000e-06|                  6.54E-08|                  6.54E-08|                           |                           |+/-6.54E-08    |Jy       |<a HREF="javascript:getReferenceInfo('2010MNRAS.408..601W','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |5.25 keV           |Broad-band measurement                                                 |                                 |Modelled datum                                           |                                        |From new raw data; NED frequency assigned to mid-point ofband in keV                                                                                               
  18|0.3-8 keV (Chandra) |          1.060000e-12|            |erg/s/cm^2^         | 1.00E+18|1.060000e-07|                          |                          |                           |                           |               |Jy       |<a HREF="javascript:getReferenceInfo('2011ApJS..192...10L','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|4.15 keV           |Broad-band measurement                                                 |03 33 36.379 -36 08 25.44 (J2000)|Flux integrated from map                                 |                                        |From reprocessed raw data; NED frequency assigned tomid-point of band in keV                                                                                       
  19|0.2-4 keV (EINSTEIN)|          1.710000e-12|            |ergs sec^-1^ cm^-2^ | 5.25E+17|3.260000e-07|                          |                          |                           |                           |               |Jy       |<a HREF="javascript:getReferenceInfo('1992ApJS...80..531F','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|2.1    keV         |Broad-band measurement; synthetic band                                 |03 31 44 -36 18 17 (B1950)       |Flux integrated from map                                 |                                        |From reprocessed raw data; Extinction-corrected for MilkyWay; NED frequency assigned to mid-point of band in keV                                                   
  20|0.5-2 keV (Swift)   |          4.000000e-13|            |erg/s/cm^2^         | 3.02E+17|1.320000e-07|                          |                          |                           |                           |               |Jy       |<a HREF="javascript:getReferenceInfo('2009ApJ...690.1322W','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|1.25 keV           |Broad-band measurement                                                 |03 33 36.4 -36 08 25.4 (J2000)   |Modelled datum                                           |                                        |From new raw data; NED frequency assigned to mid-point ofband in keV                                                                                               
  21|0.3-2 keV (XMM)     |          2.610000e-12|+/-0.03E-12 |erg/cm^2^/s         | 2.78E+17|9.390000e-07|                  1.08E-08|                  1.08E-08|                           |                           |+/-1.08E-08    |Jy       |<a HREF="javascript:getReferenceInfo('2009A&A...505..589G','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |1.15    keV        |Broad-band measurement                                                 |                                 |Modelled datum                                           |Observed flux                           |From reprocessed raw data; NED frequency assigned tomid-point of band in keV                                                                                       
  22|0.3-2 keV (Chandra) |          6.200000e-13|+/-1.3E-13  |erg/cm^2^/s         | 2.78E+17|2.230000e-07|                  4.68E-08|                  4.68E-08|                           |                           |+/-4.68E-08    |Jy       |<a HREF="javascript:getReferenceInfo('2009A&A...505..589G','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |1.15    keV        |Broad-band measurement                                                 |                                 |Modelled datum                                           |                                        |From reprocessed raw data; NED frequency assigned tomid-point of band in keV                                                                                       
  23|O VII 22.1 A (XMM)  |          2.160000e-14|+/-0.44E-14 |erg/cm^2^/s         | 1.36E+17|2.160000e+09|                  4.40E+08|                  4.40E+08|                           |                           |+/-4.40E+08    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2011ApJ...727..130K','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |22.1 A             |Line measurement; flux integrated over line; lines measured in emission|                                 |From fitting to map                                      |                                        |Averaged from previously published data                                                                                                                            
  24|NUV (GALEX) AB      |          1.200000e+01|+/-0.01     |mag                 | 1.32E+15|5.810000e-02|                  5.35E-04|                  5.35E-04|                           |                           |+/-5.35E-04    |Jy       |<a HREF="javascript:getReferenceInfo('2007ApJS..173..185G','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |2267 A             |Broad-band measurement                                                 |03 33 36.4 -36 08 25.5 (J2000)   |Total flux                                               |                                        |From new raw data                                                                                                                                                  
  25|U (Johnson)         |          1.550000e+01|+/-0.65     |milliJy             | 8.19E+14|1.550000e-02|                  6.50E-04|                  6.50E-04|                           |                           |+/-6.50E-04    |Jy       |<a HREF="javascript:getReferenceInfo('1983ApJS...52..341M','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|1 sigma                |0.366      microns |Broad-band measurement                                                 |033141.0 -361821 (B1950)         |Flux in fixed aperture                                   |29.3\" aperture                         |From new raw data                                                                                                                                                  
  26|U (Johnson)         |          9.930000e+00|+/-0.59     |milliJy             | 8.19E+14|9.930000e-03|                  5.90E-04|                  5.90E-04|                           |                           |+/-5.90E-04    |Jy       |<a HREF="javascript:getReferenceInfo('1983ApJS...52..341M','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|1 sigma                |0.366      microns |Broad-band measurement                                                 |033141.0 -361821 (B1950)         |Flux in fixed aperture                                   |22.5\" aperture                         |From new raw data                                                                                                                                                  
  27|U (U_T)             |          1.050000e+01|+/-0.08     |mag                 | 8.19E+14|1.160000e-01|                  8.45E-03|                  8.45E-03|                           |                           |+/-8.45E-03    |Jy       |<a HREF="javascript:getReferenceInfo('1991RC3.9.C...0000d','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|rms uncertainty        |3660       A       |Broad-band measurement                                                 |033142.0 -361818 (B1950)         |Multiple methods                                         |                                        |Homogenized from new and previously published data; StandardJohnson UBVRI filters assumed                                                                          
  28|U (U_T^0)           |          1.000000e+01|            |mag                 | 8.19E+14|1.780000e-01|                          |                          |                           |                           |               |Jy       |<a HREF="javascript:getReferenceInfo('1991RC3.9.C...0000d','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|3660       A       |Broad-band measurement                                                 |033142.0 -361818 (B1950)         |Multiple methods                                         |                                        |Homogenized from new and previously published data;Extinction-corrected for internal and Milky Way and K-correction applied; Standard Johnson UBVRI filters assumed
  29|B (B_T)             |          1.030000e+01|+/-0.07     |mag                 | 6.81E+14|3.170000e-01|                  2.11E-02|                  2.11E-02|                           |                           |+/-2.11E-02    |Jy       |<a HREF="javascript:getReferenceInfo('1991RC3.9.C...0000d','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|rms uncertainty        |4400       A       |Broad-band measurement                                                 |033142.0 -361818 (B1950)         |Multiple methods                                         |                                        |Homogenized from new and previously published data; StandardJohnson UBVRI filters assumed                                                                          
  30|B (Cousins) (B_26)  |          1.010000e+01|+/-0.09     |mag                 | 6.81E+14|3.790000e-01|                  3.28E-02|                  3.28E-02|                           |                           |+/-3.28E-02    |Jy       |<a HREF="javascript:getReferenceInfo('1989ESOLV.C...0000L','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|typical accuracy       |4400       A       |Broad-band measurement; photometric system transformed                 |033141 -3618.4 (B1950)           |Modelled datum                                           |See ESO-LV catalog for warning flag.    |From new raw data                                                                                                                                                  
  31|B (B_T^0)           |          9.930000e+00|            |mag                 | 6.81E+14|4.540000e-01|                          |                          |                           |                           |               |Jy       |<a HREF="javascript:getReferenceInfo('1991RC3.9.C...0000d','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|4400       A       |Broad-band measurement                                                 |033142.0 -361818 (B1950)         |Multiple methods                                         |                                        |Homogenized from new and previously published data;Extinction-corrected for internal and Milky Way and K-correction applied; Standard Johnson UBVRI filters assumed
  32|B (m_B)             |          1.020000e+01|+/-0.15     |mag                 | 6.81E+14|3.450000e-01|                  5.11E-02|                  5.11E-02|                           |                           |+/-5.11E-02    |Jy       |<a HREF="javascript:getReferenceInfo('1991RC3.9.C...0000d','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|rms uncertainty        |4400       A       |Broad-band measurement                                                 |033142.0 -361818 (B1950)         |Multiple methods                                         |                                        |Homogenized from new and previously published data; StandardJohnson UBVRI filters assumed                                                                          
  33|B (Cousins) (B_25)  |          1.020000e+01|+/-0.09     |mag                 | 6.81E+14|3.550000e-01|                  3.07E-02|                  3.07E-02|                           |                           |+/-3.07E-02    |Jy       |<a HREF="javascript:getReferenceInfo('1989ESOLV.C...0000L','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|typical accuracy       |4400       A       |Broad-band measurement; photometric system transformed                 |033141 -3618.4 (B1950)           |Modelled datum                                           |See ESO-LV catalog for warning flag.    |From new raw data                                                                                                                                                  
  34|B (Cousins) (B_T)   |          1.010000e+01|+/-0.09     |mag                 | 6.81E+14|3.970000e-01|                  3.43E-02|                  3.43E-02|                           |                           |+/-3.43E-02    |Jy       |<a HREF="javascript:getReferenceInfo('1989ESOLV.C...0000L','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|typical accuracy       |4400       A       |Broad-band measurement; photometric system transformed                 |033141 -3618.4 (B1950)           |Modelled datum                                           |See ESO-LV catalog for warning flag.    |From new raw data                                                                                                                                                  
  35|B (Johnson)         |          3.980000e+01|+/-0.79     |milliJy             | 6.69E+14|3.980000e-02|                  7.90E-04|                  7.90E-04|                           |                           |+/-7.90E-04    |Jy       |<a HREF="javascript:getReferenceInfo('1983ApJS...52..341M','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|1 sigma                |0.448      microns |Broad-band measurement                                                 |033141.0 -361821 (B1950)         |Flux in fixed aperture                                   |29.3\" aperture                         |From new raw data                                                                                                                                                  
  36|B (Johnson)         |          2.900000e+01|+/-0.62     |milliJy             | 6.69E+14|2.900000e-02|                  6.20E-04|                  6.20E-04|                           |                           |+/-6.20E-04    |Jy       |<a HREF="javascript:getReferenceInfo('1983ApJS...52..341M','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|1 sigma                |0.448      microns |Broad-band measurement                                                 |033141.0 -361821 (B1950)         |Flux in fixed aperture                                   |22.5\" aperture                         |From new raw data                                                                                                                                                  
  37|B_J                 |          1.000000e+01|            |mag                 | 6.41E+14|3.840000e-01|                          |                          |                           |                           |               |Jy       |<a HREF="javascript:getReferenceInfo('2005MNRAS.361...34D','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|4680   A           |Broad-band measurement                                                 |033335.5 -360830.4 (J2000)       |Flux in fixed aperture                                   |                                        |From new raw data                                                                                                                                                  
  38|V (Johnson)         |          9.820000e+00|            |mag                 | 5.42E+14|4.300000e-01|                          |                          |                           |                           |               |Jy       |<a HREF="javascript:getReferenceInfo('1988VIrPh.C...0000d','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|5530   A           |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                   |261.9\" aperture                        |From new raw data; Corrected for contaminating foregroundstars                                                                                                     
  39|V (Johnson)         |          4.700000e+01|+/-0.81     |milliJy             | 5.42E+14|4.700000e-02|                  8.10E-04|                  8.10E-04|                           |                           |+/-8.10E-04    |Jy       |<a HREF="javascript:getReferenceInfo('1983ApJS...52..341M','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|1 sigma                |5530   A           |Broad-band measurement                                                 |03 31 41.0 -36 18 21 (B1950)     |Flux in fixed aperture                                   |22.5\" aperture                         |From new raw data                                                                                                                                                  
  40|V (Johnson)         |          6.780000e+01|+/-1.13     |milliJy             | 5.42E+14|6.780000e-02|                  1.13E-03|                  1.13E-03|                           |                           |+/-1.13E-03    |Jy       |<a HREF="javascript:getReferenceInfo('1983ApJS...52..341M','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|1 sigma                |5530   A           |Broad-band measurement                                                 |03 31 41.0 -36 18 21 (B1950)     |Flux in fixed aperture                                   |29.3\" aperture                         |From new raw data                                                                                                                                                  
  41|V (V_T)             |          9.630000e+00|+/-0.07     |mag                 | 5.42E+14|5.120000e-01|                  3.44E-02|                  3.44E-02|                           |                           |+/-3.44E-02    |Jy       |<a HREF="javascript:getReferenceInfo('1991RC3.9.C...0000d','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|rms uncertainty        |5530       A       |Broad-band measurement                                                 |033142.0 -361818 (B1950)         |Multiple methods                                         |                                        |Homogenized from new and previously published data; StandardJohnson UBVRI filters assumed                                                                          
  42|V (LCO)             |          9.210000e+00|            |mag                 | 5.42E+14|7.540000e-01|                          |                          |                           |                           |               |Jy       |<a HREF="javascript:getReferenceInfo('2008ApJ...674..797Z','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|5530 A             |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                   |Isophotal mag                           |From new raw data; Extinction-corrected for internal andMilky Way                                                                                                  
  43|V (V_T^0)           |          9.340000e+00|            |mag                 | 5.42E+14|6.680000e-01|                          |                          |                           |                           |               |Jy       |<a HREF="javascript:getReferenceInfo('1991RC3.9.C...0000d','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|5530       A       |Broad-band measurement                                                 |033142.0 -361818 (B1950)         |Multiple methods                                         |                                        |Homogenized from new and previously published data;Extinction-corrected for internal and Milky Way and K-correction applied; Standard Johnson UBVRI filters assumed
  44|R                   |          1.020000e+01|            |mag                 | 4.68E+14|2.640000e-01|                          |                          |                           |                           |               |Jy       |<a HREF="javascript:getReferenceInfo('2005MNRAS.361...34D','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|6400   A           |Broad-band measurement                                                 |033335.5 -360830.4 (J2000)       |Flux in fixed aperture                                   |                                        |From new raw data                                                                                                                                                  
  45|R (Cousins) (R_T)   |          8.790000e+00|+/-0.09     |mag                 | 4.68E+14|9.400000e-01|                  8.12E-02|                  8.12E-02|                           |                           |+/-8.12E-02    |Jy       |<a HREF="javascript:getReferenceInfo('1989ESOLV.C...0000L','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|typical accuracy       |6400       A       |Broad-band measurement; photometric system transformed                 |033141 -3618.4 (B1950)           |Modelled datum                                           |See ESO-LV catalog for warning flag.    |From new raw data                                                                                                                                                  
  48|R' (Johnson)        |          9.340000e+00|            |mag                 | 4.48E+14|5.110000e-01|                          |                          |                           |                           |               |Jy       |<a HREF="javascript:getReferenceInfo('1988VIrPh.C...0000d','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|6690   A           |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                   |261.9\" aperture                        |From new raw data; Corrected for contaminating foregroundstars                                                                                                     
  49|R (Johnson)         |          8.470000e+01|+/-2.17     |milliJy             | 4.28E+14|8.470000e-02|                  2.17E-03|                  2.17E-03|                           |                           |+/-2.17E-03    |Jy       |<a HREF="javascript:getReferenceInfo('1983ApJS...52..341M','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|1 sigma                |7000   A           |Broad-band measurement                                                 |03 31 41.0 -36 18 21 (B1950)     |Flux in fixed aperture                                   |22.5\" aperture                         |From new raw data                                                                                                                                                  
  50|R (Johnson)         |          1.230000e+02|+/-3.16     |milliJy             | 4.28E+14|1.230000e-01|                  3.16E-03|                  3.16E-03|                           |                           |+/-3.16E-03    |Jy       |<a HREF="javascript:getReferenceInfo('1983ApJS...52..341M','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|1 sigma                |7000   A           |Broad-band measurement                                                 |03 31 41.0 -36 18 21 (B1950)     |Flux in fixed aperture                                   |29.3\" aperture                         |From new raw data                                                                                                                                                  
  52|I_t_                |          8.350000e+00|            |mag                 | 3.80E+14|1.090000e+00|                          |                          |                           |                           |               |Jy       |<a HREF="javascript:getReferenceInfo('1997AJ....113...22G','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|8060       A       |Broad-band measurement                                                 |033141.8 -361824. (B1950)        |Total flux                                               |                                        |Averaged new and previously published data; Corrected forcontaminating foreground stars                                                                            
  53|I_corr_             |          8.240000e+00|+/-0.11     |mag                 | 3.80E+14|1.200000e+00|                  5.03E-01|                  5.03E-01|                           |                           |+/-5.03E-01    |Jy       |<a HREF="javascript:getReferenceInfo('1997AJ....113...22G','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |8060       A       |Broad-band measurement                                                 |033141.8 -361824. (B1950)        |Total flux                                               |                                        |Averaged new and previously published data;Extinction-corrected for internal and Milky Way and K-correction applied                                                
  54|I                   |          9.730000e+00|            |mag                 | 3.79E+14|3.270000e-01|                          |                          |                           |                           |               |Jy       |<a HREF="javascript:getReferenceInfo('2005MNRAS.361...34D','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|7900   A           |Broad-band measurement                                                 |033335.5 -360830.4 (J2000)       |Flux in fixed aperture                                   |                                        |From new raw data                                                                                                                                                  
  55|I                   |          8.320000e+00|            |mag                 | 3.79E+14|1.200000e+00|                          |                          |                           |                           |               |Jy       |<a HREF="javascript:getReferenceInfo('2007ApJS..172..599S','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|7900 A             |Broad-band measurement                                                 |03 33 36.3 -36 08 23 (J2000)     |Total flux                                               |                                        |Averaged new and previously published data;Extinction-corrected for Milky Way; Standard Cousins R_C, I_C filters assumed                                           
  56|I                   |          8.420000e+00|+/-0.04     |mag                 | 3.79E+14|1.090000e+00|                  4.03E-02|                  4.03E-02|                           |                           |+/-4.03E-02    |Jy       |<a HREF="javascript:getReferenceInfo('2007ApJS..172..599S','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |7900 A             |Broad-band measurement                                                 |03 33 36.3 -36 08 23 (J2000)     |Total flux                                               |Observed magnitude                      |Averaged new and previously published data; Standard CousinsR_C, I_C filters assumed                                                                               
  57|I (LCO)             |          8.050000e+00|            |mag                 | 3.79E+14|1.540000e+00|                          |                          |                           |                           |               |Jy       |<a HREF="javascript:getReferenceInfo('2008ApJ...674..797Z','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|7900 A             |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                   |Isophotal mag                           |From new raw data; Extinction-corrected for internal andMilky Way                                                                                                  
  58|I' (Johnson)        |          8.850000e+00|            |mag                 | 3.75E+14|6.460000e-01|                          |                          |                           |                           |               |Jy       |<a HREF="javascript:getReferenceInfo('1988VIrPh.C...0000d','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|8000   A           |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                   |261.9\" aperture                        |From new raw data; Corrected for contaminating foregroundstars                                                                                                     
  59|I (KPNO)            |          8.320000e+00|+/-0.06     |mag                 | 3.65E+14|1.200000e+00|                  6.62E-02|                  6.62E-02|                           |                           |+/-6.62E-02    |Jy       |<a HREF="javascript:getReferenceInfo('2006ApJ...653..969T','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |8204.53   A        |Broad-band measurement                                                 |                                 |Total flux                                               |                                        |Averaged new and previously published data;Extinction-corrected for internal and Milky Way                                                                         
  60|I (Johnson)         |          1.250000e+02|+/-4.12     |milliJy             | 3.33E+14|1.250000e-01|                  4.12E-03|                  4.12E-03|                           |                           |+/-4.12E-03    |Jy       |<a HREF="javascript:getReferenceInfo('1983ApJS...52..341M','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|1 sigma                |9000   A           |Broad-band measurement                                                 |03 31 41.0 -36 18 21 (B1950)     |Flux in fixed aperture                                   |22.5\" aperture                         |From new raw data                                                                                                                                                  
  61|I (Johnson)         |          1.670000e+02|+/-5.38     |milliJy             | 3.33E+14|1.670000e-01|                  5.38E-03|                  5.38E-03|                           |                           |+/-5.38E-03    |Jy       |<a HREF="javascript:getReferenceInfo('1983ApJS...52..341M','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|1 sigma                |9000   A           |Broad-band measurement                                                 |03 31 41.0 -36 18 21 (B1950)     |Flux in fixed aperture                                   |29.3\" aperture                         |From new raw data                                                                                                                                                  
  62|J (ESO/SPM)         |          1.490000e+02|+/-9.89     |milliJy             | 2.50E+14|1.490000e-01|                  9.89E-03|                  9.89E-03|                           |                           |+/-9.89E-03    |Jy       |<a HREF="javascript:getReferenceInfo('1995ApJ...453..616S','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|rms uncertainty        |1.198      microns |Broad-band measurement                                                 |033141.9 -361824 (B1950)         |Flux in fixed aperture                                   |15\" aperture                           |From new raw data                                                                                                                                                  
  63|J (RGO)             |          9.220000e+00|+/-0.09     |mag                 | 2.50E+14|3.360000e-01|                  2.91E-02|                  2.91E-02|                           |                           |+/-2.91E-02    |Jy       |<a HREF="javascript:getReferenceInfo('1973MNRAS.164..155G','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |1.2 microns        |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                   |37.8\" aperture                         |From new raw data                                                                                                                                                  
  64|J                   |          9.100000e+00|+/-0.12     |mag                 | 2.50E+14|3.760000e-01|                  4.39E-02|                  4.39E-02|                           |                           |+/-4.39E-02    |Jy       |<a HREF="javascript:getReferenceInfo('1976MNRAS.175..191G','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |1.2     microns    |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                   |25\" aperture                           |From new raw data; Extinction-corrected for Milky Way;derived from a flux in a different band and a color                                                          
  65|J (RGO)             |          8.950000e+00|+/-0.09     |mag                 | 2.50E+14|4.310000e-01|                  3.73E-02|                  3.73E-02|                           |                           |+/-3.73E-02    |Jy       |<a HREF="javascript:getReferenceInfo('1973MNRAS.164..155G','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |1.2 microns        |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                   |37.8\" aperture                         |From new raw data                                                                                                                                                  
  66|J (RGO)             |          1.060000e+01|+/-0.10     |mag                 | 2.50E+14|9.530000e-02|                  9.19E-03|                  9.19E-03|                           |                           |+/-9.19E-03    |Jy       |<a HREF="javascript:getReferenceInfo('1973MNRAS.164..155G','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |1.2 microns        |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                   |12\" aperture;Low quality data          |From new raw data                                                                                                                                                  
  69|J (Johnson)         |          8.750000e+00|+/-0.03     |mag                 | 2.42E+14|5.070000e-01|                  1.42E-02|                  1.42E-02|                           |                           |+/-1.42E-02    |Jy       |<a HREF="javascript:getReferenceInfo('1977HarvU.T00M....A','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |1.24    microns    |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                   |55.8\" aperture                         |From new raw data; derived from a flux in a different bandand a color                                                                                              
  70|J (Johnson)         |          9.330000e+00|+/-0.03     |mag                 | 2.42E+14|2.970000e-01|                  8.32E-03|                  8.32E-03|                           |                           |+/-8.32E-03    |Jy       |<a HREF="javascript:getReferenceInfo('1977HarvU.T00M....A','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |1.24    microns    |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                   |28.6\" aperture                         |From new raw data; derived from a flux in a different bandand a color                                                                                              
  73|J_tot (2MASS LGA)   |          7.360000e+00|+/-0.026    |mag                 | 2.40E+14|1.810000e+00|                  4.38E-02|                  4.38E-02|                           |                           |+/-4.38E-02    |Jy       |<a HREF="javascript:getReferenceInfo('2003AJ....125..525J','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|1 sigma uncert.        |1.25      microns  |Broad-band measurement                                                 |033336.46 -360826.4 (J2000)      |Total flux                                               |                                        |From new raw data                                                                                                                                                  
  75|J (Johnson)         |          3.220000e+02|+/-8.4      |milliJy             | 2.38E+14|3.220000e-01|                  8.40E-03|                  8.40E-03|                           |                           |+/-8.40E-03    |Jy       |<a HREF="javascript:getReferenceInfo('1983ApJS...52..341M','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|1 sigma                |1.26    microns    |Broad-band measurement                                                 |03 31 41.0 -36 18 21 (B1950)     |Flux in fixed aperture                                   |22.8\" aperture                         |From new raw data                                                                                                                                                  
  76|J (Johnson)         |          2.570000e+02|+/-6.8      |milliJy             | 2.38E+14|2.570000e-01|                  6.80E-03|                  6.80E-03|                           |                           |+/-6.80E-03    |Jy       |<a HREF="javascript:getReferenceInfo('1983ApJS...52..341M','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|1 sigma                |1.26    microns    |Broad-band measurement                                                 |03 31 41.0 -36 18 21 (B1950)     |Flux in fixed aperture                                   |13.7\" aperture                         |From new raw data                                                                                                                                                  
  77|J (Johnson)         |          1.860000e+02|+/-5.0      |milliJy             | 2.38E+14|1.860000e-01|                  5.00E-03|                  5.00E-03|                           |                           |+/-5.00E-03    |Jy       |<a HREF="javascript:getReferenceInfo('1983ApJS...52..341M','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|1 sigma                |1.26    microns    |Broad-band measurement                                                 |03 31 41.0 -36 18 21 (B1950)     |Flux in fixed aperture                                   |9.1\" aperture                          |From new raw data                                                                                                                                                  
  78|H (ESO/SPM)         |          2.490000e+02|+/-16.59    |milliJy             | 1.90E+14|2.490000e-01|                  1.66E-02|                  1.66E-02|                           |                           |+/-1.66E-02    |Jy       |<a HREF="javascript:getReferenceInfo('1995ApJ...453..616S','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|rms uncertainty        |1.580      microns |Broad-band measurement                                                 |033141.9 -361824 (B1950)         |Flux in fixed aperture                                   |15\" aperture                           |From new raw data                                                                                                                                                  
  79|H (Johnson)         |          4.390000e+02|+/-11.1     |milliJy             | 1.87E+14|4.390000e-01|                  1.11E-02|                  1.11E-02|                           |                           |+/-1.11E-02    |Jy       |<a HREF="javascript:getReferenceInfo('1983ApJS...52..341M','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|1 sigma                |1.60    microns    |Broad-band measurement                                                 |03 31 41.0 -36 18 21 (B1950)     |Flux in fixed aperture                                   |13.7\" aperture                         |From new raw data                                                                                                                                                  
  80|H (Johnson)         |          5.350000e+02|+/-15.1     |milliJy             | 1.87E+14|5.340000e-01|                  1.51E-02|                  1.51E-02|                           |                           |+/-1.51E-02    |Jy       |<a HREF="javascript:getReferenceInfo('1983ApJS...52..341M','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|1 sigma                |1.60    microns    |Broad-band measurement                                                 |03 31 41.0 -36 18 21 (B1950)     |Flux in fixed aperture                                   |22.8\" aperture                         |From new raw data                                                                                                                                                  
  81|H (Johnson)         |          3.200000e+02|+/-8.1      |milliJy             | 1.87E+14|3.200000e-01|                  8.10E-03|                  8.10E-03|                           |                           |+/-8.10E-03    |Jy       |<a HREF="javascript:getReferenceInfo('1983ApJS...52..341M','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|1 sigma                |1.60    microns    |Broad-band measurement                                                 |03 31 41.0 -36 18 21 (B1950)     |Flux in fixed aperture                                   |9.1\" aperture                          |From new raw data                                                                                                                                                  
  82|H                   |          8.190000e+00|+/-0.12     |mag                 | 1.83E+14|5.460000e-01|                  6.38E-02|                  6.38E-02|                           |                           |+/-6.38E-02    |Jy       |<a HREF="javascript:getReferenceInfo('1976MNRAS.175..191G','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |1.64    microns    |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                   |25\" aperture                           |From new raw data; Extinction-corrected for Milky Way;derived from a flux in a different band and a color                                                          
  83|H (RGO)             |          8.220000e+00|+/-0.09     |mag                 | 1.83E+14|5.310000e-01|                  4.59E-02|                  4.59E-02|                           |                           |+/-4.59E-02    |Jy       |<a HREF="javascript:getReferenceInfo('1973MNRAS.164..155G','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |1.64 microns       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                   |37.8\" aperture                         |From new raw data                                                                                                                                                  
  84|H (RGO)             |          9.590000e+00|+/-0.14     |mag                 | 1.83E+14|1.500000e-01|                  2.07E-02|                  2.07E-02|                           |                           |+/-2.07E-02    |Jy       |<a HREF="javascript:getReferenceInfo('1973MNRAS.164..155G','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |1.64 microns       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                   |12\" aperture;Low quality data          |From new raw data                                                                                                                                                  
  85|H (RGO)             |          8.210000e+00|+/-0.08     |mag                 | 1.83E+14|5.360000e-01|                  4.10E-02|                  4.10E-02|                           |                           |+/-4.10E-02    |Jy       |<a HREF="javascript:getReferenceInfo('1973MNRAS.164..155G','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |1.64 microns       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                   |37.8\" aperture                         |From new raw data                                                                                                                                                  
  88|H_tot (2MASS LGA)   |          6.740000e+00|+/-0.031    |mag                 | 1.82E+14|2.070000e+00|                  5.99E-02|                  5.99E-02|                           |                           |+/-5.99E-02    |Jy       |<a HREF="javascript:getReferenceInfo('2003AJ....125..525J','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|1 sigma uncert.        |1.65      microns  |Broad-band measurement                                                 |033336.46 -360826.4 (J2000)      |Total flux                                               |                                        |From new raw data                                                                                                                                                  
  90|H (HCO)             |          7.510000e+00|+/-0.03     |mag                 | 1.82E+14|9.710000e-01|                  2.72E-02|                  2.72E-02|                           |                           |+/-2.72E-02    |Jy       |<a HREF="javascript:getReferenceInfo('1981MNRAS.195p...1A','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |1.65    microns    |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                   |110.0\" aperture                        |From new raw data                                                                                                                                                  
  91|H (HCO)             |          7.190000e+00|+/-0.03     |mag                 | 1.82E+14|1.300000e+00|                  3.65E-02|                  3.65E-02|                           |                           |+/-3.65E-02    |Jy       |<a HREF="javascript:getReferenceInfo('1981MNRAS.195p...1A','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |1.65    microns    |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                   |165.2\" aperture                        |From new raw data                                                                                                                                                  
  92|H (HCO)             |          7.470000e+00|+/-0.03     |mag                 | 1.82E+14|1.010000e+00|                  2.82E-02|                  2.82E-02|                           |                           |+/-2.82E-02    |Jy       |<a HREF="javascript:getReferenceInfo('1981MNRAS.195p...1A','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |1.65    microns    |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                   |110.6\" aperture                        |From new raw data                                                                                                                                                  
  93|H (HCO)             |          7.680000e+00|+/-0.03     |mag                 | 1.82E+14|8.300000e-01|                  2.33E-02|                  2.33E-02|                           |                           |+/-2.33E-02    |Jy       |<a HREF="javascript:getReferenceInfo('1981MNRAS.195p...1A','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |1.65    microns    |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                   |83.6\" aperture                         |From new raw data                                                                                                                                                  
  94|H (HCO)             |          8.010000e+00|+/-0.03     |mag                 | 1.82E+14|6.130000e-01|                  1.72E-02|                  1.72E-02|                           |                           |+/-1.72E-02    |Jy       |<a HREF="javascript:getReferenceInfo('1981MNRAS.195p...1A','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |1.65    microns    |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                   |50.4\" aperture                         |From new raw data                                                                                                                                                  
  95|H (HCO)             |          7.940000e+00|+/-0.03     |mag                 | 1.82E+14|6.540000e-01|                  1.83E-02|                  1.83E-02|                           |                           |+/-1.83E-02    |Jy       |<a HREF="javascript:getReferenceInfo('1981MNRAS.195p...1A','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |1.65    microns    |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                   |55.8\" aperture                         |Transformed from previously published data                                                                                                                         
  96|H (Johnson)         |          8.450000e+00|+/-0.03     |mag                 | 1.82E+14|4.480000e-01|                  1.26E-02|                  1.26E-02|                           |                           |+/-1.26E-02    |Jy       |<a HREF="javascript:getReferenceInfo('1977HarvU.T00M....A','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |1.65    microns    |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                   |28.6\" aperture                         |From new raw data; derived from a flux in a different bandand a color                                                                                              
  97|H (Johnson)         |          7.940000e+00|+/-0.03     |mag                 | 1.82E+14|7.170000e-01|                  2.01E-02|                  2.01E-02|                           |                           |+/-2.01E-02    |Jy       |<a HREF="javascript:getReferenceInfo('1977HarvU.T00M....A','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |1.65    microns    |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                   |55.8\" aperture                         |From new raw data; derived from a flux in a different bandand a color                                                                                              
 100|H_2 1-0 S(1) (VLT)  |                      |<0.78E-18   |W m^-2^             | 1.41E+14|            |                          |                          |                    7.8E+07|                           |<7.80E+07      |Jy       |<a HREF="javascript:getReferenceInfo('2005ApJ...633..105D','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|2.1218   microns   |Line measurement; flux integrated over line; lines measured in emission|03 33 36.4 -36 08 25 (J2000)     |Flux in fixed aperture                                   |Flux extracted in 1\" length of 1\" slit|From new raw data                                                                                                                                                  
 101|K (VLT/ISAAC)       |          9.800000e+00|            |mag                 | 1.39E+14|8.020000e-02|                          |                          |                           |                           |               |Jy       |<a HREF="javascript:getReferenceInfo('2005ApJ...633..105D','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|2.16   microns     |Broad-band measurement                                                 |03 33 36.4 -36 08 25 (J2000)     |Flux in fixed aperture                                   |Mag extracted in 1\" length of 1\" slit |From new raw data                                                                                                                                                  
 106|K_tot (2MASS LGA)   |          6.370000e+00|+/-0.036    |mag                 | 1.38E+14|1.880000e+00|                  6.35E-02|                  6.35E-02|                           |                           |+/-6.35E-02    |Jy       |<a HREF="javascript:getReferenceInfo('2003AJ....125..525J','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|1 sigma uncert.        |2.17      microns  |Broad-band measurement                                                 |033336.46 -360826.4 (J2000)      |Total flux                                               |                                        |From new raw data                                                                                                                                                  
 108|K (RGO)             |          7.710000e+00|+/-0.09     |mag                 | 1.37E+14|5.360000e-01|                  4.63E-02|                  4.63E-02|                           |                           |+/-4.63E-02    |Jy       |<a HREF="javascript:getReferenceInfo('1973MNRAS.164..155G','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |2.19 microns       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                   |37.8\" aperture                         |From new raw data                                                                                                                                                  
 109|K                   |          7.750000e+00|+/-0.12     |mag                 | 1.37E+14|5.160000e-01|                  6.03E-02|                  6.03E-02|                           |                           |+/-6.03E-02    |Jy       |<a HREF="javascript:getReferenceInfo('1976MNRAS.175..191G','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |2.19    microns    |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                   |25\" aperture                           |From new raw data; Extinction-corrected for Milky Way                                                                                                              
 110|K (RGO)             |          7.810000e+00|+/-0.09     |mag                 | 1.37E+14|4.890000e-01|                  4.22E-02|                  4.22E-02|                           |                           |+/-4.22E-02    |Jy       |<a HREF="javascript:getReferenceInfo('1973MNRAS.164..155G','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |2.19 microns       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                   |37.8\" aperture                         |From new raw data                                                                                                                                                  
 111|K (RGO)             |          8.880000e+00|+/-0.08     |mag                 | 1.37E+14|1.820000e-01|                  1.39E-02|                  1.39E-02|                           |                           |+/-1.39E-02    |Jy       |<a HREF="javascript:getReferenceInfo('1973MNRAS.164..155G','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |2.19 microns       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                   |12\" aperture                           |From new raw data                                                                                                                                                  
 112|K (ESO/SPM)         |          2.640000e+02|+/-17.59    |milliJy             | 1.36E+14|2.640000e-01|                  1.76E-02|                  1.76E-02|                           |                           |+/-1.76E-02    |Jy       |<a HREF="javascript:getReferenceInfo('1995ApJ...453..616S','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|rms uncertainty        |2.210      microns |Broad-band measurement                                                 |033141.9 -361824 (B1950)         |Flux in fixed aperture                                   |15\" aperture                           |From new raw data                                                                                                                                                  
 113|K (Johnson)         |          7.990000e+00|+/-0.03     |mag                 | 1.35E+14|4.250000e-01|                  1.19E-02|                  1.19E-02|                           |                           |+/-1.19E-02    |Jy       |<a HREF="javascript:getReferenceInfo('1977HarvU.T00M....A','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |2.22    microns    |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                   |28.6\" aperture                         |From new raw data                                                                                                                                                  
 114|K (Johnson)         |          3.250000e+02|+/-5.7      |milliJy             | 1.35E+14|3.250000e-01|                  5.70E-03|                  5.70E-03|                           |                           |+/-5.70E-03    |Jy       |<a HREF="javascript:getReferenceInfo('1983ApJS...52..341M','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|1 sigma                |2.22    microns    |Broad-band measurement                                                 |03 31 41.0 -36 18 21 (B1950)     |Flux in fixed aperture                                   |9.1\" aperture                          |From new raw data                                                                                                                                                  
 115|K (Johnson)         |          4.260000e+02|+/-7.3      |milliJy             | 1.35E+14|4.260000e-01|                  7.30E-03|                  7.30E-03|                           |                           |+/-7.30E-03    |Jy       |<a HREF="javascript:getReferenceInfo('1983ApJS...52..341M','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|1 sigma                |2.22    microns    |Broad-band measurement                                                 |03 31 41.0 -36 18 21 (B1950)     |Flux in fixed aperture                                   |13.7\" aperture                         |From new raw data                                                                                                                                                  
 116|K (Johnson)         |          4.790000e+02|+/-9.4      |milliJy             | 1.35E+14|4.790000e-01|                  9.40E-03|                  9.40E-03|                           |                           |+/-9.40E-03    |Jy       |<a HREF="javascript:getReferenceInfo('1983ApJS...52..341M','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|1 sigma                |2.22    microns    |Broad-band measurement                                                 |03 31 41.0 -36 18 21 (B1950)     |Flux in fixed aperture                                   |22.8\" aperture                         |From new raw data                                                                                                                                                  
 117|K (Johnson)         |          7.580000e+00|+/-0.03     |mag                 | 1.35E+14|6.200000e-01|                  1.74E-02|                  1.74E-02|                           |                           |+/-1.74E-02    |Jy       |<a HREF="javascript:getReferenceInfo('1977HarvU.T00M....A','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |2.22    microns    |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                   |55.8\" aperture                         |From new raw data                                                                                                                                                  
 118|L                   |          6.280000e+00|+/-0.12     |mag                 | 8.82E+13|8.610000e-01|                  1.01E-01|                  1.01E-01|                           |                           |+/-1.01E-01    |Jy       |<a HREF="javascript:getReferenceInfo('1976MNRAS.175..191G','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |3.4     microns    |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                   |25\" aperture                           |From new raw data; Extinction-corrected for Milky Way;derived from a flux in a different band and a color                                                          
 119|L (RGO)             |          6.750000e+00|+/-0.74     |mag                 | 8.57E+13|5.590000e-01|                  5.46E-01|                  5.46E-01|                           |                           |+/-5.46E-01    |Jy       |<a HREF="javascript:getReferenceInfo('1973MNRAS.164..155G','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |3.5 microns        |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                   |37.8\" aperture                         |From new raw data                                                                                                                                                  
 120|L (RGO)             |          6.230000e+00|+/-0.25     |mag                 | 8.57E+13|9.020000e-01|                  2.34E-01|                  2.34E-01|                           |                           |+/-2.34E-01    |Jy       |<a HREF="javascript:getReferenceInfo('1973MNRAS.164..155G','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |3.5 microns        |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                   |37.8\" aperture                         |From new raw data                                                                                                                                                  
 121|L (RGO)             |          7.460000e+00|+/-0.18     |mag                 | 8.57E+13|2.910000e-01|                  5.24E-02|                  5.24E-02|                           |                           |+/-5.24E-02    |Jy       |<a HREF="javascript:getReferenceInfo('1973MNRAS.164..155G','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |3.5 microns        |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                   |12\" aperture                           |From new raw data                                                                                                                                                  
 122|L (Johnson)         |          3.240000e+02|+/-5.9      |milliJy             | 8.47E+13|3.240000e-01|                  5.90E-03|                  5.90E-03|                           |                           |+/-5.90E-03    |Jy       |<a HREF="javascript:getReferenceInfo('1983ApJS...52..341M','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|1 sigma                |3.54    microns    |Broad-band measurement                                                 |03 31 41.0 -36 18 21 (B1950)     |Flux in fixed aperture                                   |13.7\" aperture                         |From new raw data                                                                                                                                                  
 123|L (Johnson)         |          2.550000e+02|+/-5.8      |milliJy             | 8.47E+13|2.550000e-01|                  5.80E-03|                  5.80E-03|                           |                           |+/-5.80E-03    |Jy       |<a HREF="javascript:getReferenceInfo('1983ApJS...52..341M','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|1 sigma                |3.54    microns    |Broad-band measurement                                                 |03 31 41.0 -36 18 21 (B1950)     |Flux in fixed aperture                                   |9.1\" aperture                          |From new raw data                                                                                                                                                  
 124|L (Johnson)         |          4.340000e+02|+/-10.3     |milliJy             | 8.47E+13|4.340000e-01|                  1.03E-02|                  1.03E-02|                           |                           |+/-1.03E-02    |Jy       |<a HREF="javascript:getReferenceInfo('1983ApJS...52..341M','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|1 sigma                |3.54    microns    |Broad-band measurement                                                 |03 31 41.0 -36 18 21 (B1950)     |Flux in fixed aperture                                   |22.8\" aperture                         |From new raw data                                                                                                                                                  
 125|3.6 microns (IRAC)  |          7.230000e+00|+/-0.07     |mag                 | 8.44E+13|3.600000e-01|                  2.32E-02|                  2.32E-02|                           |                           |+/-2.32E-02    |Jy       |<a HREF="javascript:getReferenceInfo('2010ApJS..187..172G','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |3.550 microns      |Broad-band measurement                                                 |03 33 36.39 -36 08 25.8 (J2000)  |Flux in fixed aperture                                   |                                        |From new raw data                                                                                                                                                  
 126|4.5 microns (IRAC)  |          6.850000e+00|+/-0.06     |mag                 | 6.67E+13|3.270000e-01|                  1.81E-02|                  1.81E-02|                           |                           |+/-1.81E-02    |Jy       |<a HREF="javascript:getReferenceInfo('2010ApJS..187..172G','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |4.493 microns      |Broad-band measurement                                                 |03 33 36.39 -36 08 25.8 (J2000)  |Flux in fixed aperture                                   |                                        |From new raw data                                                                                                                                                  
 127|M (Johnson)         |          2.920000e+02|+/-28.6     |milliJy             | 6.25E+13|2.920000e-01|                  2.86E-02|                  2.86E-02|                           |                           |+/-2.86E-02    |Jy       |<a HREF="javascript:getReferenceInfo('1983ApJS...52..341M','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|1 sigma                |4.8     microns    |Broad-band measurement                                                 |03 31 41.0 -36 18 21 (B1950)     |Flux in fixed aperture                                   |9.1\" aperture                          |From new raw data                                                                                                                                                  
 128|5.5 microns (IRS)   |          7.290000e-01|+/-1.26E-01 |Jy                  | 5.45E+13|7.290000e-01|                  1.26E-01|                  1.26E-01|                           |                           |+/-1.26E-01    |Jy       |<a HREF="javascript:getReferenceInfo('2009ApJ...705...14D','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |5.5 microns        |Broad-band measurement                                                 |                                 |Flux integrated from map                                 |                                        |From reprocessed raw data                                                                                                                                          
 129|5.8 microns (IRAC)  |          5.700000e+00|+/-0.08     |mag                 | 5.23E+13|6.040000e-01|                  4.45E-02|                  4.45E-02|                           |                           |+/-4.45E-02    |Jy       |<a HREF="javascript:getReferenceInfo('2010ApJS..187..172G','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |5.731 microns      |Broad-band measurement                                                 |03 33 36.39 -36 08 25.8 (J2000)  |Flux in fixed aperture                                   |                                        |From new raw data                                                                                                                                                  
 130|6 microns (IRS)     |          3.200000e-01|            |Jy                  | 5.00E+13|3.200000e-01|                          |                          |                           |                           |               |Jy       |<a HREF="javascript:getReferenceInfo('2006ApJ...653.1129B','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|6   microns        |Broad-band measurement                                                 |03 33 36.37 -36 08 25.5 (J2000)  |Flux integrated from map                                 |                                        |From new raw data                                                                                                                                                  
 131|6 microns (ISO)     |                      |<0.5582     |Jy                  | 5.00E+13|            |                          |                          |                    5.6E-01|                           |<5.58E-01      |Jy       |<a HREF="javascript:getReferenceInfo('2004A&A...418..465L','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|3 sigma                |6   microns        |Broad-band measurement                                                 |                                 |Flux integrated from map                                 |                                        |From reprocessed raw data                                                                                                                                          
 132|PAH 6.2 microns IRS |          2.740000e-19|+/-10  %    |W cm^-2^            | 4.84E+13|2.740000e+11|                  2.74E+10|                  2.74E+10|                           |                           |+/-2.74E+10    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2006ApJ...653.1129B','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|estimated error        |6.2   microns      |Line measurement; flux integrated over line                            |03 33 36.37 -36 08 25.5 (J2000)  |Flux integrated from map                                 |                                        |From new raw data                                                                                                                                                  
 133|PAH 6.2 (Spitzer)   |          1.730000e-18|+/-1E-20    |W/cm^2^             | 4.84E+13|1.730000e+09|                  1.00E+07|                  1.00E+07|                           |                           |+/-1.00E+07    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2009ApJ...701..658W','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |6.2 microns        |Line measurement; flux integrated over line; lines measured in emission|03 33 36.4 -36 08 25 (J2000)     |Flux in fixed aperture                                   |                                        |From reprocessed raw data                                                                                                                                          
 134|6.2 microns (IRS)   |          3.730000e-14|+/-180E-17  |W/m^2^              | 4.84E+13|3.730000e+12|                  1.80E+11|                  1.80E+11|                           |                           |+/-1.80E+11    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2010ApJS..187..172G','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|1 sigma                |6.2 microns        |Line measurement; flux integrated over line; lines measured in emission|03 33 36.39 -36 08 25.8 (J2000)  |Flux integrated from map                                 |                                        |From new raw data                                                                                                                                                  
 135|PAH 6.2 (Spitzer)   |          4.230000e-19|+/-0.56E-20 |W/cm^2^             | 4.84E+13|4.230000e+11|                  5.60E+09|                  5.60E+09|                           |                           |+/-5.60E+09    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2011ApJ...728...45L','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |6.2 microns        |Line measurement; flux integrated over line; lines measured in emission|                                 |Flux integrated from map                                 |                                        |From reprocessed raw data                                                                                                                                          
 136|7 microns (ISOCAM)  |          3.690000e+03|+/-616.6    |milliJy             | 4.44E+13|3.690000e+00|                  6.17E-01|                  6.17E-01|                           |                           |+/-6.17E-01    |Jy       |<a HREF="javascript:getReferenceInfo('2001A&A...369..473R','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |7.0        microns |Broad-band measurement                                                 |                                 |Flux integrated from map                                 |                                        |From new raw data                                                                                                                                                  
 138|7.4 microns (IRS)   |          4.330000e-14|+/-580E-17  |W/m^2^              | 4.05E+13|4.330000e+12|                  5.80E+11|                  5.80E+11|                           |                           |+/-5.80E+11    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2010ApJS..187..172G','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|1 sigma                |7.4 microns        |Line measurement; flux integrated over line; lines measured in emission|03 33 36.39 -36 08 25.8 (J2000)  |Flux integrated from map                                 |                                        |From new raw data                                                                                                                                                  
 139|7.6 microns (IRS)   |          4.890000e-14|+/-260E-17  |W/m^2^              | 3.94E+13|4.890000e+12|                  2.60E+11|                  2.60E+11|                           |                           |+/-2.60E+11    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2010ApJS..187..172G','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|1 sigma                |7.6 microns        |Line measurement; flux integrated over line; lines measured in emission|03 33 36.39 -36 08 25.8 (J2000)  |Flux integrated from map                                 |                                        |From new raw data                                                                                                                                                  
 140|PAH 7.7 microns IRS |          6.370000e-19|+/-10  %    |W cm^-2^            | 3.89E+13|6.370000e+11|                  6.37E+10|                  6.37E+10|                           |                           |+/-6.37E+10    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2006ApJ...653.1129B','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|estimated error        |7.7   microns      |Line measurement; flux integrated over line                            |03 33 36.37 -36 08 25.5 (J2000)  |Flux integrated from map                                 |                                        |From new raw data                                                                                                                                                  
 141|PAH 7.7 (Spitzer)   |          1.350000e-18|+/-2.54E-20 |W/cm^2^             | 3.89E+13|1.350000e+12|                  2.54E+10|                  2.54E+10|                           |                           |+/-2.54E+10    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2011ApJ...728...45L','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |7.7 microns        |Line measurement; flux integrated over line; lines measured in emission|                                 |Flux integrated from map                                 |                                        |From reprocessed raw data                                                                                                                                          
 142|7.8 microns         |                      |+/-32  %    |W cm^-2^ micron ^-1^| 3.84E+13|1.400000e+00|                  4.49E-01|                  4.49E-01|                           |                           |+/-4.49E-01    |Jy       |<a HREF="javascript:getReferenceInfo('1982ApJ...260...70F','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |7.8     microns    |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                   |12.6\" aperture                         |From new raw data; measurement modified from published value                                                                                                       
 143|7.8 microns (IRS)   |          5.610000e-14|+/-310E-17  |W/m^2^              | 3.84E+13|5.610000e+12|                  3.10E+11|                  3.10E+11|                           |                           |+/-3.10E+11    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2010ApJS..187..172G','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|1 sigma                |7.8 microns        |Line measurement; flux integrated over line; lines measured in emission|03 33 36.39 -36 08 25.8 (J2000)  |Flux integrated from map                                 |                                        |From new raw data                                                                                                                                                  
 144|8.0 microns (IRAC)  |          3.250000e+00|+/-0.09     |mag                 | 3.81E+13|3.210000e+00|                  2.66E-01|                  2.66E-01|                           |                           |+/-2.66E-01    |Jy       |<a HREF="javascript:getReferenceInfo('2010ApJS..187..172G','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |7.872 microns      |Broad-band measurement                                                 |03 33 36.39 -36 08 25.8 (J2000)  |Flux in fixed aperture                                   |                                        |From new raw data                                                                                                                                                  
 145|8.3 microns (IRS)   |          1.720000e-14|+/-190E-17  |W/m^2^              | 3.61E+13|1.720000e+12|                  1.90E+11|                  1.90E+11|                           |                           |+/-1.90E+11    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2010ApJS..187..172G','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|1 sigma                |8.3 microns        |Line measurement; flux integrated over line; lines measured in emission|03 33 36.39 -36 08 25.8 (J2000)  |Flux integrated from map                                 |                                        |From new raw data                                                                                                                                                  
 146|8.6 microns TIMMI2  |          4.000000e-01|+/-10  %    |Jy                  | 3.49E+13|4.000000e-01|                  4.00E-02|                  4.00E-02|                           |                           |+/-4.00E-02    |Jy       |<a HREF="javascript:getReferenceInfo('2004A&A...414..123S','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |8.6   microns      |Broad-band measurement                                                 |                                 |From multi-aperture data                                 |                                        |From new raw data                                                                                                                                                  
 147|PAH 8.6 microns IRS |          1.300000e-19|+/-10  %    |W cm^-2^            | 3.49E+13|1.300000e+11|                  1.30E+10|                  1.30E+10|                           |                           |+/-1.30E+10    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2006ApJ...653.1129B','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|estimated error        |8.6   microns      |Line measurement; flux integrated over line                            |03 33 36.37 -36 08 25.5 (J2000)  |Flux integrated from map                                 |                                        |From new raw data                                                                                                                                                  
 148|8.6 microns (IRS)   |          2.440000e-14|+/-84E-17   |W/m^2^              | 3.49E+13|2.440000e+12|                  8.40E+10|                  8.40E+10|                           |                           |+/-8.40E+10    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2010ApJS..187..172G','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|1 sigma                |8.6 microns        |Line measurement; flux integrated over line; lines measured in emission|03 33 36.39 -36 08 25.8 (J2000)  |Flux integrated from map                                 |                                        |From new raw data                                                                                                                                                  
 149|PAH 8.6 (Spitzer)   |          3.660000e-19|+/-1.13E-20 |W/cm^2^             | 3.49E+13|3.660000e+11|                  1.13E+10|                  1.13E+10|                           |                           |+/-1.13E+10    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2011ApJ...728...45L','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |8.6 microns        |Line measurement; flux integrated over line; lines measured in emission|                                 |Flux integrated from map                                 |                                        |From reprocessed raw data                                                                                                                                          
 150|8.6 microns         |                      |+/-12  %    |W cm^-2^ micron ^-1^| 3.49E+13|1.050000e+00|                  1.26E-01|                  1.26E-01|                           |                           |+/-1.26E-01    |Jy       |<a HREF="javascript:getReferenceInfo('1982ApJ...260...70F','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |8.6     microns    |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                   |12.6\" aperture                         |From new raw data; measurement modified from published value                                                                                                       
 151|8.9 microns (TIMMI2)|          4.100000e+02|+/-82       |milliJy             | 3.43E+13|4.100000e-01|                  8.20E-02|                  8.20E-02|                           |                           |+/-8.20E-02    |Jy       |<a HREF="javascript:getReferenceInfo('2005A&A...438..803G','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |8.73   microns     |Broad-band measurement                                                 |03 33 36.4 -36 08 25 (J2000)     |Flux in fixed aperture                                   |                                        |From new raw data                                                                                                                                                  
 152|9.6 microns         |                      |+/-14  %    |W cm^-2^ micron ^-1^| 3.12E+13|5.990000e-01|                  8.39E-02|                  8.39E-02|                           |                           |+/-8.39E-02    |Jy       |<a HREF="javascript:getReferenceInfo('1982ApJ...260...70F','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |9.6     microns    |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                   |12.6\" aperture                         |From new raw data; measurement modified from published value                                                                                                       
 153|10 microns (IRS)    |          1.230000e+00|+/-7.41E-02 |Jy                  | 3.00E+13|1.230000e+00|                  7.41E-02|                  7.41E-02|                           |                           |+/-7.41E-02    |Jy       |<a HREF="javascript:getReferenceInfo('2009ApJ...705...14D','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |10 microns         |Broad-band measurement                                                 |                                 |Flux integrated from map                                 |                                        |From reprocessed raw data                                                                                                                                          
 154|10.4 microns TIMMI2 |          4.400000e+02|+/-88       |milliJy             | 2.89E+13|4.400000e-01|                  8.80E-02|                  8.80E-02|                           |                           |+/-8.80E-02    |Jy       |<a HREF="javascript:getReferenceInfo('2005A&A...438..803G','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |10.38   microns    |Broad-band measurement                                                 |03 33 36.4 -36 08 25 (J2000)     |Flux in fixed aperture                                   |                                        |From new raw data                                                                                                                                                  
 155|N (CTIO)            |          3.210000e+02|+/-15  %    |milliJy             | 2.89E+13|3.210000e-01|                  4.82E-02|                  4.82E-02|                           |                           |+/-4.82E-02    |Jy       |<a HREF="javascript:getReferenceInfo('2009ApJ...702.1127R','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|estimated error        |10.36 microns      |Broad-band measurement                                                 |                                 |From fitting to map                                      |Nuclear flux                            |From new raw data                                                                                                                                                  
 156|10.4 microns        |                      |+/-9   %    |W cm^-2^ micron ^-1^| 2.88E+13|9.710000e-01|                  8.74E-02|                  8.74E-02|                           |                           |+/-8.74E-02    |Jy       |<a HREF="javascript:getReferenceInfo('1982ApJ...260...70F','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |10.4     microns   |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                   |12.6\" aperture                         |From new raw data; measurement modified from published value                                                                                                       
 157|10.4 microns TIMMI2 |          4.600000e-01|+/-10  %    |Jy                  | 2.88E+13|4.600000e-01|                  4.60E-02|                  4.60E-02|                           |                           |+/-4.60E-02    |Jy       |<a HREF="javascript:getReferenceInfo('2004A&A...414..123S','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |10.4   microns     |Broad-band measurement                                                 |                                 |From multi-aperture data                                 |                                        |From new raw data                                                                                                                                                  
 158|[S IV] 10.51 (IRS)  |          1.860000e-13|+/-0.78E-14 |erg/s/cm^2^         | 2.85E+13|1.860000e+10|                  7.80E+08|                  7.80E+08|                           |                           |+/-7.80E+08    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2010ApJ...709.1257T','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |10.51 microns      |Line measurement; flux integrated over line; lines measured in emission|03 33 36.4 -36 08 25 (J2000)     |Flux integrated from map                                 |SH module                               |From new raw data                                                                                                                                                  
 159|[S IV] (TIMMI2)     |                      |<1.7E-20    |W cm^-2^            | 2.85E+13|            |                          |                          |                    1.7E+10|                           |<1.70E+10      |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2004A&A...414..123S','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|3 sigma                |10.511   microns   |Line measurement; flux integrated over line                            |                                 |Flux integrated from map                                 |3\" aperture                            |From new raw data                                                                                                                                                  
 160|[S IV] (ISO)        |          2.600000e-20|            |W cm^-2^            | 2.85E+13|2.600000e+10|                          |                          |                           |                           |               |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2004A&A...414..123S','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|10.511   microns   |Line measurement; flux integrated over line                            |                                 |Flux integrated from map                                 |14\"x20\" aper; from 2002A&A...393..821S|Averaged from previously published data                                                                                                                            
 161|10 microns          |                      |+/-8   %    |W cm^-2^ micron ^-1^| 2.83E+13|8.980000e-01|                  7.18E-02|                  7.18E-02|                           |                           |+/-7.18E-02    |Jy       |<a HREF="javascript:getReferenceInfo('1982ApJ...260...70F','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |10.6     microns   |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                   |12.6\" aperture                         |From new raw data; measurement modified from published value                                                                                                       
 162|PAH 11.2 (Spitzer)  |          1.200000e-18|+/-3E-20    |W/cm^2^             | 2.68E+13|1.200000e+09|                  3.00E+07|                  3.00E+07|                           |                           |+/-3.00E+07    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2009ApJ...701..658W','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |11.2 microns       |Line measurement; flux integrated over line; lines measured in emission|03 33 36.4 -36 08 25 (J2000)     |Flux in fixed aperture                                   |                                        |From reprocessed raw data                                                                                                                                          
 163|11.2 microns (IRS)  |          8.390000e-15|+/-42E-17   |W/m^2^              | 2.68E+13|8.390000e+11|                  4.20E+10|                  4.20E+10|                           |                           |+/-4.20E+10    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2010ApJS..187..172G','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|1 sigma                |11.2 microns       |Line measurement; flux integrated over line; lines measured in emission|03 33 36.39 -36 08 25.8 (J2000)  |Flux integrated from map                                 |                                        |From new raw data                                                                                                                                                  
 164|PAH2 (VLT)          |          4.230000e+02|+/-7.8      |milliJy             | 2.66E+13|4.230000e-01|                  7.80E-03|                  7.80E-03|                           |                           |+/-7.80E-03    |Jy       |<a HREF="javascript:getReferenceInfo('2014MNRAS.439.1648A','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |11.25   microns    |Broad-band measurement                                                 |053.401667 -36.140278 (J2000)    |Flux in fixed aperture                                   |Nuclear flux                            |From reprocessed raw data                                                                                                                                          
 165|11.3 microns (ISO)  |          1.250000e-18|            |W cm^-2^            | 2.65E+13|1.250000e+12|                          |                          |                           |                           |               |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2004A&A...414..123S','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|11.3   microns     |Line measurement; flux integrated over line                            |                                 |Flux integrated from map                                 |24\" aperture                           |Averaged from previously published data                                                                                                                            
 166|11.3 microns TIMMI2 |                      |<11E-20     |W cm^-2^            | 2.65E+13|            |                          |                          |                    1.1E+11|                           |<1.10E+11      |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2004A&A...414..123S','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|11.3   microns     |Line measurement; flux integrated over line                            |                                 |Flux integrated from map                                 |3\" slit                                |From new raw data                                                                                                                                                  
 167|11.3 microns (IRS)  |          2.510000e-14|+/-110E-17  |W/m^2^              | 2.65E+13|2.510000e+12|                  1.10E+11|                  1.10E+11|                           |                           |+/-1.10E+11    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2010ApJS..187..172G','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|1 sigma                |11.3 microns       |Line measurement; flux integrated over line; lines measured in emission|03 33 36.39 -36 08 25.8 (J2000)  |Flux integrated from map                                 |                                        |From new raw data                                                                                                                                                  
 168|PAH 11.3 (Spitzer)  |          7.030000e-19|+/-1.5E-20  |W/cm^2^             | 2.65E+13|7.030000e+11|                  1.50E+10|                  1.50E+10|                           |                           |+/-1.50E+10    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2011ApJ...728...45L','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |11.3 microns       |Line measurement; flux integrated over line; lines measured in emission|                                 |Flux integrated from map                                 |                                        |From reprocessed raw data                                                                                                                                          
 169|PAH 11.3 microns IRS|          4.600000e-19|+/-10  %    |W cm^-2^            | 2.65E+13|4.600000e+11|                  4.60E+10|                  4.60E+10|                           |                           |+/-4.60E+10    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2006ApJ...653.1129B','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|estimated error        |11.3   microns     |Line measurement; flux integrated over line                            |03 33 36.37 -36 08 25.5 (J2000)  |Flux integrated from map                                 |                                        |From new raw data                                                                                                                                                  
 170|11.4 microns        |                      |+/-12  %    |W cm^-2^ micron ^-1^| 2.63E+13|9.710000e-01|                  1.17E-01|                  1.17E-01|                           |                           |+/-1.17E-01    |Jy       |<a HREF="javascript:getReferenceInfo('1982ApJ...260...70F','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |11.4     microns   |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                   |12.6\" aperture                         |From new raw data; measurement modified from published value                                                                                                       
 171|11.9 microns TIMMI2 |          5.100000e+02|+/-102      |milliJy             | 2.57E+13|5.100000e-01|                  1.02E-01|                  1.02E-01|                           |                           |+/-1.02E-01    |Jy       |<a HREF="javascript:getReferenceInfo('2005A&A...438..803G','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |11.66   microns    |Broad-band measurement                                                 |03 33 36.4 -36 08 25 (J2000)     |Flux in fixed aperture                                   |                                        |From new raw data                                                                                                                                                  
 172|11.9 microns TIMMI2 |          6.060000e+02|+/-15  %    |milliJy             | 2.52E+13|6.060000e-01|                  9.09E-02|                  9.09E-02|                           |                           |+/-9.09E-02    |Jy       |<a HREF="javascript:getReferenceInfo('2008A&A...484..341R','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|estimated error        |11.9 microns       |Broad-band measurement                                                 |03 33 36.4 -36 08 25.5 (J2000)   |Flux in fixed aperture                                   |                                        |From new raw data                                                                                                                                                  
 173|12 microns (VLTI)   |          5.100000e-01|            |Jy                  | 2.50E+13|5.100000e-01|                          |                          |                           |                           |               |Jy       |<a HREF="javascript:getReferenceInfo('2009A&A...502...67T','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|12 microns         |Broad-band measurement                                                 |03 33 36.38 -36 08 25.7 (J2000)  |Total flux                                               |                                        |From new raw data                                                                                                                                                  
 174|12.0 microns (IRS)  |          1.240000e-14|+/-64E-17   |W/m^2^              | 2.50E+13|1.240000e+12|                  6.40E+10|                  6.40E+10|                           |                           |+/-6.40E+10    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2010ApJS..187..172G','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|1 sigma                |12.0 microns       |Line measurement; flux integrated over line; lines measured in emission|03 33 36.39 -36 08 25.8 (J2000)  |Flux integrated from map                                 |                                        |From new raw data                                                                                                                                                  
 175|12 microns (IRAS)   |          5.120000e+00|+/-0.031    |Jy                  | 2.50E+13|5.120000e+00|                  3.10E-02|                  3.10E-02|                           |                           |+/-3.10E-02    |Jy       |<a HREF="javascript:getReferenceInfo('2003AJ....126.1607S','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|1 sigma                |12   microns       |Broad-band measurement                                                 |03 33 36.5 -36 08 23 (J2000)     |Total flux                                               |Size, Method, Flag codes: RZ;see paper  |From reprocessed raw data                                                                                                                                          
 178|NEII_1 (VLT)        |          4.910000e+02|+/-27.0     |milliJy             | 2.44E+13|4.910000e-01|                  2.70E-02|                  2.70E-02|                           |                           |+/-2.70E-02    |Jy       |<a HREF="javascript:getReferenceInfo('2014MNRAS.439.1648A','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |12.27   microns    |Broad-band measurement                                                 |053.401667 -36.140278 (J2000)    |Flux in fixed aperture                                   |Nuclear flux                            |From reprocessed raw data                                                                                                                                          
 179|12.9 microns TIMMI2 |          1.100000e+02|+/-220      |milliJy             | 2.43E+13|1.100000e-01|                  2.20E-01|                  2.20E-01|                           |                           |+/-2.20E-01    |Jy       |<a HREF="javascript:getReferenceInfo('2005A&A...438..803G','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |12.35   microns    |Broad-band measurement                                                 |03 33 36.4 -36 08 25 (J2000)     |Flux in fixed aperture                                   |                                        |From new raw data                                                                                                                                                  
 180|12.4 microns        |                      |+/-18  %    |W cm^-2^ micron ^-1^| 2.42E+13|1.410000e+00|                  2.54E-01|                  2.54E-01|                           |                           |+/-2.54E-01    |Jy       |<a HREF="javascript:getReferenceInfo('1982ApJ...260...70F','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |12.4     microns   |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                   |12.6\" aperture                         |From new raw data; measurement modified from published value                                                                                                       
 181|12.6 microns (IRS)  |          2.590000e-14|+/-180E-17  |W/m^2^              | 2.38E+13|2.590000e+12|                  1.80E+11|                  1.80E+11|                           |                           |+/-1.80E+11    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2010ApJS..187..172G','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|1 sigma                |12.6 microns       |Line measurement; flux integrated over line; lines measured in emission|03 33 36.39 -36 08 25.8 (J2000)  |Flux integrated from map                                 |                                        |From new raw data                                                                                                                                                  
 182|[Ne II] 12.81 (IRS) |          1.400000e-19|+/-3.27E-21 |W/cm^2^             | 2.34E+13|1.400000e+11|                  3.27E+09|                  3.27E+09|                           |                           |+/-3.27E+09    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2009ApJS..184..230B','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |12.81 microns      |Line measurement; flux integrated over line; lines measured in emission|03 33 36.37 -36 08 25.5 (J2000)  |Flux integrated from map                                 |                                        |From new raw data                                                                                                                                                  
 183|[Ne II] (TIMMI2)    |                      |<1.8E-20    |W cm^-2^            | 2.34E+13|            |                          |                          |                    1.8E+10|                           |<1.80E+10      |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2004A&A...414..123S','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|3 sigma                |12.814   microns   |Line measurement; flux integrated over line                            |                                 |Flux integrated from map                                 |3\" aperture                            |From new raw data                                                                                                                                                  
 184|[Ne II] (ISO)       |          4.090000e-19|            |W cm^-2^            | 2.34E+13|4.090000e+11|                          |                          |                           |                           |               |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2004A&A...414..123S','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|12.814   microns   |Line measurement; flux integrated over line                            |                                 |Flux integrated from map                                 |14\"x27\" aper; from 2002A&A...393..821S|Averaged from previously published data                                                                                                                            
 185|[Ne II] 12.81 (IRS) |          1.430000e-12|+/-3.79E-14 |erg/s/cm^2^         | 2.34E+13|1.430000e+11|                  3.79E+09|                  3.79E+09|                           |                           |+/-3.79E+09    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2010ApJ...709.1257T','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |12.81 microns      |Line measurement; flux integrated over line; lines measured in emission|03 33 36.4 -36 08 25 (J2000)     |Flux integrated from map                                 |SH module                               |From new raw data                                                                                                                                                  
 186|[Ne II] 12.81 (IRS) |          1.620000e-19|+/-17.48E-21|W/cm^2^             | 2.34E+13|1.620000e+11|                  1.75E+10|                  1.75E+10|                           |                           |+/-1.75E+10    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2010ApJ...716.1151W','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|1 sigma                |12.81 microns      |Line measurement; flux integrated over line; lines measured in emission|                                 |Flux integrated from map                                 |                                        |From reprocessed raw data                                                                                                                                          
 187|[Ne II] 12.8 Spitzer|          1.560000e-12|            |erg/cm^2^/s         | 2.34E+13|1.560000e+11|                          |                          |                           |                           |               |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2010ApJ...725.2270P','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|12.81 microns      |Line measurement; flux integrated over line; lines measured in emission|03 33 36.4 -36 08 25 (J2000)     |From fitting to map                                      |                                        |From reprocessed raw data                                                                                                                                          
 188|[Ne II] 12.81       |          1.400000e-19|            |W/cm^2^             | 2.34E+13|1.400000e+11|                          |                          |                           |                           |               |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2011ApJS..195...17W','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|12.81 microns      |Line measurement; flux integrated over line; lines measured in emission|                                 |Not reported in paper                                    |                                        |Averaged from previously published data                                                                                                                            
 189|NEII (VLT)          |          5.980000e+02|+/-16.7     |milliJy             | 2.34E+13|5.980000e-01|                  1.67E-02|                  1.67E-02|                           |                           |+/-1.67E-02    |Jy       |<a HREF="javascript:getReferenceInfo('2014MNRAS.439.1648A','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |12.81   microns    |Broad-band measurement                                                 |053.401667 -36.140278 (J2000)    |Flux in fixed aperture                                   |Nuclear flux                            |From reprocessed raw data                                                                                                                                          
 190|NEII (VLT)          |          6.400000e+02|+/-20.3     |milliJy             | 2.34E+13|6.400000e-01|                  2.03E-02|                  2.03E-02|                           |                           |+/-2.03E-02    |Jy       |<a HREF="javascript:getReferenceInfo('2014MNRAS.439.1648A','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |12.81   microns    |Broad-band measurement                                                 |053.401667 -36.140278 (J2000)    |Flux in fixed aperture                                   |Nuclear flux                            |From reprocessed raw data                                                                                                                                          
 191|NEII_2 (VLT)        |          5.020000e+02|+/-11.1     |milliJy             | 2.30E+13|5.020000e-01|                  1.11E-02|                  1.11E-02|                           |                           |+/-1.11E-02    |Jy       |<a HREF="javascript:getReferenceInfo('2014MNRAS.439.1648A','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |13.04   microns    |Broad-band measurement                                                 |053.401667 -36.140278 (J2000)    |Flux in fixed aperture                                   |Nuclear flux                            |From reprocessed raw data                                                                                                                                          
 192|PAH 14.2 microns IRS|          6.200000e-20|+/-10  %    |W cm^-2^            | 2.11E+13|6.200000e+10|                  6.20E+09|                  6.20E+09|                           |                           |+/-6.20E+09    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2006ApJ...653.1129B','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|estimated error        |14.2   microns     |Line measurement; flux integrated over line                            |03 33 36.37 -36 08 25.5 (J2000)  |Flux integrated from map                                 |                                        |From new raw data                                                                                                                                                  
 193|[Ne V] 14.3 Spitzer |          2.160000e-16|+/-10.5E-18 |W/m^2^              | 2.10E+13|2.160000e+10|                  1.05E+09|                  1.05E+09|                           |                           |+/-1.05E+09    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2011ApJ...730...28P','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |14.3 microns       |Line measurement; flux integrated over line; lines measured in emission|53.4015 -36.1404 (J2000)         |Flux integrated from map                                 |                                        |From new raw data                                                                                                                                                  
 194|[Ne V] 14.32        |          2.200000e-20|+/-0.06E-20 |W/cm^2^             | 2.09E+13|2.200000e+10|                  6.00E+08|                  6.00E+08|                           |                           |+/-6.00E+08    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2007ApJ...664...71D','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|statistical error      |14.32   microns    |Line measurement; flux integrated over line; lines measured in emission|                                 |Flux integrated from map                                 |                                        |From reprocessed raw data                                                                                                                                          
 195|[Ne V] 14.32 (IRS)  |          1.910000e-13|+/-0.61E-14 |erg/s/cm^2^         | 2.09E+13|1.910000e+10|                  6.10E+08|                  6.10E+08|                           |                           |+/-6.10E+08    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2010ApJ...709.1257T','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |14.32 microns      |Line measurement; flux integrated over line; lines measured in emission|03 33 36.4 -36 08 25 (J2000)     |Flux integrated from map                                 |SH module                               |From new raw data                                                                                                                                                  
 196|[Ne V] 14.32 (IRS)  |          2.240000e-20|+/-1.97E-21 |W/cm^2^             | 2.09E+13|2.240000e+10|                  1.97E+09|                  1.97E+09|                           |                           |+/-1.97E+09    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2010ApJ...716.1151W','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|1 sigma                |14.32 microns      |Line measurement; flux integrated over line; lines measured in emission|                                 |Flux integrated from map                                 |                                        |From reprocessed raw data                                                                                                                                          
 197|[Ne V] 14.3 Spitzer |          1.900000e-13|            |erg/cm^2^/s         | 2.09E+13|1.900000e+10|                          |                          |                           |                           |               |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2010ApJ...725.2270P','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|14.32 microns      |Line measurement; flux integrated over line; lines measured in emission|03 33 36.4 -36 08 25 (J2000)     |From fitting to map                                      |                                        |From reprocessed raw data                                                                                                                                          
 198|[Ne V] 14.32        |          1.880000e-20|            |W/cm^2^             | 2.09E+13|1.880000e+10|                          |                          |                           |                           |               |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2011ApJS..195...17W','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|14.32 microns      |Line measurement; flux integrated over line; lines measured in emission|                                 |Not reported in paper                                    |                                        |Averaged from previously published data                                                                                                                            
 199|14.7 microns (IRS)  |          2.690000e+00|+/-1.28E-01 |Jy                  | 2.04E+13|2.690000e+00|                  1.28E-01|                  1.28E-01|                           |                           |+/-1.28E-01    |Jy       |<a HREF="javascript:getReferenceInfo('2009ApJ...705...14D','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |14.7 microns       |Broad-band measurement                                                 |                                 |Flux integrated from map                                 |                                        |From reprocessed raw data                                                                                                                                          
 200|LW3 (ISOCAM)        |          3.100000e+03|+/-20       |milliJy             | 2.00E+13|3.100000e+00|                  6.21E-01|                  6.21E-01|                           |                           |+/-6.21E-01    |Jy       |<a HREF="javascript:getReferenceInfo('2004A&A...419..501F','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|estimated error        |15.0   microns     |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                   |40.0\" diameter aperture                |From reprocessed raw data                                                                                                                                          
 201|15 microns (ISO)    |          4.440000e+03|+/-764.5    |milliJy             | 2.00E+13|4.440000e+00|                  7.65E-01|                  7.65E-01|                           |                           |+/-7.65E-01    |Jy       |<a HREF="javascript:getReferenceInfo('2001A&A...369..473R','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |15.0       microns |Broad-band measurement                                                 |                                 |Flux integrated from map                                 |                                        |From new raw data                                                                                                                                                  
 202|15 microns (IRS)    |          1.550000e+00|            |Jy                  | 2.00E+13|1.550000e+00|                          |                          |                           |                           |               |Jy       |<a HREF="javascript:getReferenceInfo('2006ApJ...653.1129B','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|15   microns       |Broad-band measurement                                                 |03 33 36.37 -36 08 25.5 (J2000)  |Flux integrated from map                                 |                                        |From new raw data                                                                                                                                                  
 203|[Ne III] 15.56 (IRS)|          6.130000e-13|+/-0.51E-14 |erg/s/cm^2^         | 1.93E+13|6.130000e+10|                  5.10E+08|                  5.10E+08|                           |                           |+/-5.10E+08    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2010ApJ...709.1257T','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |15.56 microns      |Line measurement; flux integrated over line; lines measured in emission|03 33 36.4 -36 08 25 (J2000)     |Flux integrated from map                                 |SH module                               |From new raw data                                                                                                                                                  
 204|[Ne III] 15.56 (IRS)|          6.110000e-20|+/-0.90E-21 |W/cm^2^             | 1.93E+13|6.110000e+10|                  9.00E+08|                  9.00E+08|                           |                           |+/-9.00E+08    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2010ApJ...716.1151W','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|1 sigma                |15.56 microns      |Line measurement; flux integrated over line; lines measured in emission|                                 |Flux integrated from map                                 |                                        |From reprocessed raw data                                                                                                                                          
 205|[Ne III] 15.5 (IRS) |          5.950000e-20|+/-0.92E-21 |W/cm^2^             | 1.93E+13|5.950000e+10|                  9.20E+08|                  9.20E+08|                           |                           |+/-9.20E+08    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2009ApJS..184..230B','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |15.55 microns      |Line measurement; flux integrated over line; lines measured in emission|03 33 36.37 -36 08 25.5 (J2000)  |Flux integrated from map                                 |                                        |From new raw data                                                                                                                                                  
 206|[NeIII] 15.6 Spitzer|          6.100000e-13|            |erg/cm^2^/s         | 1.93E+13|6.100000e+10|                          |                          |                           |                           |               |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2010ApJ...725.2270P','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|15.56 microns      |Line measurement; flux integrated over line; lines measured in emission|03 33 36.4 -36 08 25 (J2000)     |From fitting to map                                      |                                        |From reprocessed raw data                                                                                                                                          
 207|[Ne III] 15.56      |          5.950000e-20|            |W/cm^2^             | 1.93E+13|5.950000e+10|                          |                          |                           |                           |               |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2011ApJS..195...17W','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|15.56 microns      |Line measurement; flux integrated over line; lines measured in emission|                                 |Not reported in paper                                    |                                        |Averaged from previously published data                                                                                                                            
 208|17.0 microns (IRS)  |          1.220000e-14|+/-82E-17   |W/m^2^              | 1.76E+13|1.220000e+12|                  8.20E+10|                  8.20E+10|                           |                           |+/-8.20E+10    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2010ApJS..187..172G','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|1 sigma                |17.0 microns       |Line measurement; flux integrated over line; lines measured in emission|03 33 36.39 -36 08 25.8 (J2000)  |Flux integrated from map                                 |                                        |From new raw data                                                                                                                                                  
 209|PAH 17 microns IRS  |          5.590000e-19|+/-10  %    |W cm^-2^            | 1.76E+13|5.590000e+11|                  5.59E+10|                  5.59E+10|                           |                           |+/-5.59E+10    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2006ApJ...653.1129B','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|estimated error        |17   microns       |Line measurement; flux integrated over line                            |03 33 36.37 -36 08 25.5 (J2000)  |Flux integrated from map                                 |                                        |From new raw data                                                                                                                                                  
 210|Qa (GeminiS)        |          6.400000e+02|+/-25  %    |milliJy             | 1.64E+13|6.400000e-01|                  1.60E-01|                  1.60E-01|                           |                           |+/-1.60E-01    |Jy       |<a HREF="javascript:getReferenceInfo('2009ApJ...702.1127R','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|estimated error        |18.33 microns      |Broad-band measurement                                                 |                                 |From fitting to map                                      |Nuclear flux                            |From new raw data                                                                                                                                                  
 211|[S III] 18.71 (IRS) |          5.120000e-13|+/-0.57E-14 |erg/s/cm^2^         | 1.60E+13|5.120000e+10|                  5.70E+08|                  5.70E+08|                           |                           |+/-5.70E+08    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2010ApJ...709.1257T','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |18.71 microns      |Line measurement; flux integrated over line; lines measured in emission|03 33 36.4 -36 08 25 (J2000)     |Flux integrated from map                                 |SH module                               |From new raw data                                                                                                                                                  
 212|[S III] 18.71 (IRS) |          5.370000e-20|+/-3.58E-21 |W/cm^2^             | 1.60E+13|5.370000e+10|                  3.58E+09|                  3.58E+09|                           |                           |+/-3.58E+09    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2009ApJS..184..230B','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |18.71 microns      |Line measurement; flux integrated over line; lines measured in emission|03 33 36.37 -36 08 25.5 (J2000)  |Flux integrated from map                                 |                                        |From new raw data                                                                                                                                                  
 213|[S III] 18.71       |          5.730000e-20|+/-0.05E-20 |W/cm^2^             | 1.60E+13|5.730000e+10|                  5.00E+08|                  5.00E+08|                           |                           |+/-5.00E+08    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2007ApJ...664...71D','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|statistical error      |18.71   microns    |Line measurement; flux integrated over line; lines measured in emission|                                 |Flux integrated from map                                 |                                        |From reprocessed raw data                                                                                                                                          
 214|20 microns (IRS)    |          4.890000e+00|+/-1.18E-01 |Jy                  | 1.50E+13|4.890000e+00|                  1.18E-01|                  1.18E-01|                           |                           |+/-1.18E-01    |Jy       |<a HREF="javascript:getReferenceInfo('2009ApJ...705...14D','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |20 microns         |Broad-band measurement                                                 |                                 |Flux integrated from map                                 |                                        |From reprocessed raw data                                                                                                                                          
 215|20 microns          |                      |+/-60  %    |W cm^-2^ micron ^-1^| 1.50E+13|1.600000e+00|                  9.63E-01|                  9.63E-01|                           |                           |+/-9.63E-01    |Jy       |<a HREF="javascript:getReferenceInfo('1982ApJ...260...70F','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |20       microns   |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                   |12.6\" aperture                         |From new raw data; measurement modified from published value                                                                                                       
 216|[Ne V] 24.32        |          5.360000e-20|+/-0.06E-20 |W/cm^2^             | 1.23E+13|5.360000e+10|                  6.00E+08|                  6.00E+08|                           |                           |+/-6.00E+08    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2007ApJ...664...71D','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|statistical error      |24.31   microns    |Line measurement; flux integrated over line; lines measured in emission|                                 |Flux integrated from map                                 |                                        |From reprocessed raw data                                                                                                                                          
 217|[Ne V] 24.32 (IRS)  |          9.750000e-13|+/-13.2E-14 |erg/s/cm^2^         | 1.23E+13|9.750000e+10|                  1.32E+10|                  1.32E+10|                           |                           |+/-1.32E+10    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2010ApJ...709.1257T','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |24.32 microns      |Line measurement; flux integrated over line; lines measured in emission|03 33 36.4 -36 08 25 (J2000)     |Flux integrated from map                                 |LH module                               |From new raw data                                                                                                                                                  
 218|[Ne V] 24.32 (IRS)  |          3.850000e-20|+/-1.50E-21 |W/cm^2^             | 1.23E+13|2.240000e+10|                  1.50E+09|                  1.50E+09|                           |                           |+/-1.50E+09    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2010ApJ...716.1151W','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|1 sigma                |24.32 microns      |Line measurement; flux integrated over line; lines measured in emission|                                 |Flux integrated from map                                 |                                        |From reprocessed raw data                                                                                                                                          
 220|25 microns (IRAS)   |          1.430000e+01|+/-0.038    |Jy                  | 1.20E+13|1.430000e+01|                  3.80E-02|                  3.80E-02|                           |                           |+/-3.80E-02    |Jy       |<a HREF="javascript:getReferenceInfo('2003AJ....126.1607S','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|1 sigma                |25   microns       |Broad-band measurement                                                 |03 33 36.5 -36 08 23 (J2000)     |Total flux                                               |Size, Method, Flag codes: RZ;see paper  |From reprocessed raw data                                                                                                                                          
 223|[O IV] 25.89 (IRS)  |          3.650000e-12|+/-26.9E-14 |erg/s/cm^2^         | 1.16E+13|3.650000e+11|                  2.69E+10|                  2.69E+10|                           |                           |+/-2.69E+10    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2010ApJ...709.1257T','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |25.89 microns      |Line measurement; flux integrated over line; lines measured in emission|03 33 36.4 -36 08 25 (J2000)     |Flux integrated from map                                 |LH module                               |From new raw data                                                                                                                                                  
 224|[O IV] 25.89 (IRS)  |          1.450000e-19|+/-8.89E-21 |W/cm^2^             | 1.16E+13|1.450000e+11|                  8.89E+09|                  8.89E+09|                           |                           |+/-8.89E+09    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2010ApJ...716.1151W','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|1 sigma                |25.89 microns      |Line measurement; flux integrated over line; lines measured in emission|                                 |Flux integrated from map                                 |                                        |From reprocessed raw data                                                                                                                                          
 225|[O IV] 25.9 Spitzer |          1.510000e-12|            |erg/cm^2^/s         | 1.16E+13|1.510000e+11|                          |                          |                           |                           |               |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2010ApJ...725.2270P','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|25.89 microns      |Line measurement; flux integrated over line; lines measured in emission|03 33 36.4 -36 08 25 (J2000)     |From fitting to map                                      |                                        |From reprocessed raw data                                                                                                                                          
 226|[O IV] 25.89 Spitzer|          1.580000e-12|+/-0.12e-12 |erg/cm^2^/s         | 1.16E+13|1.580000e+11|                  1.20E+10|                  1.20E+10|                           |                           |+/-1.20E+10    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2009ApJ...698..623D','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |25.89 microns      |Line measurement; flux integrated over line; lines measured in emission|                                 |Flux integrated from map                                 |                                        |From reprocessed raw data                                                                                                                                          
 227|[O IV] 25.89        |          1.420000e-19|            |W/cm^2^             | 1.16E+13|1.420000e+11|                          |                          |                           |                           |               |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2011ApJS..195...17W','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|25.89 microns      |Line measurement; flux integrated over line; lines measured in emission|                                 |Not reported in paper                                    |                                        |Averaged from previously published data                                                                                                                            
 228|[Fe II] 25.99       |          2.220000e-20|            |W/cm^2^             | 1.15E+13|2.220000e+10|                          |                          |                           |                           |               |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2011ApJS..195...17W','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|25.99 microns      |Line measurement; flux integrated over line; lines measured in emission|                                 |Not reported in paper                                    |                                        |Averaged from previously published data                                                                                                                            
 229|30 microns (IRS)    |          1.230000e+01|+/-3.43E-01 |Jy                  | 9.99E+12|1.230000e+01|                  3.43E-01|                  3.43E-01|                           |                           |+/-3.43E-01    |Jy       |<a HREF="javascript:getReferenceInfo('2009ApJ...705...14D','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |30 microns         |Broad-band measurement                                                 |                                 |Flux integrated from map                                 |                                        |From reprocessed raw data                                                                                                                                          
 230|30 microns (IRS)    |          9.610000e+00|            |Jy                  | 9.99E+12|9.610000e+00|                          |                          |                           |                           |               |Jy       |<a HREF="javascript:getReferenceInfo('2006ApJ...653.1129B','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|30   microns       |Broad-band measurement                                                 |03 33 36.37 -36 08 25.5 (J2000)  |Flux integrated from map                                 |                                        |From new raw data                                                                                                                                                  
 231|[S III] 33.48 (IRS) |          7.200000e-12|+/-102.E-14 |erg/s/cm^2^         | 8.95E+12|7.200000e+11|                  1.02E+11|                  1.02E+11|                           |                           |+/-1.02E+11    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2010ApJ...709.1257T','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |33.48 microns      |Line measurement; flux integrated over line; lines measured in emission|03 33 36.4 -36 08 25 (J2000)     |Flux integrated from map                                 |LH module                               |From new raw data                                                                                                                                                  
 232|[S III] 33.48       |          2.720000e-19|+/-0.38E-20 |W/cm^2^             | 8.95E+12|2.720000e+11|                  3.80E+09|                  3.80E+09|                           |                           |+/-3.80E+09    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2007ApJ...664...71D','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|statistical error      |33.48   microns    |Line measurement; flux integrated over line; lines measured in emission|                                 |Flux integrated from map                                 |                                        |From reprocessed raw data                                                                                                                                          
 233|[S III] 33.48       |          2.470000e-19|            |W/cm^2^             | 8.95E+12|2.470000e+11|                          |                          |                           |                           |               |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2011ApJS..195...17W','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|33.48 microns      |Line measurement; flux integrated over line; lines measured in emission|                                 |Not reported in paper                                    |                                        |Averaged from previously published data                                                                                                                            
 234|[S III] 33.48 (IRS) |          2.470000e-19|+/-12.17E-21|W/cm^2^             | 8.95E+12|2.470000e+11|                  1.22E+10|                  1.22E+10|                           |                           |+/-1.22E+10    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2009ApJS..184..230B','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |33.48 microns      |Line measurement; flux integrated over line; lines measured in emission|03 33 36.37 -36 08 25.5 (J2000)  |Flux integrated from map                                 |                                        |From new raw data                                                                                                                                                  
 235|[Si II] 34.28       |          5.000000e-19|            |W/cm^2^             | 8.75E+12|5.000000e+11|                          |                          |                           |                           |               |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2011ApJS..195...17W','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|34.28 microns      |Line measurement; flux integrated over line; lines measured in emission|                                 |Not reported in paper                                    |                                        |Averaged from previously published data                                                                                                                            
 236|[Si II] 34.82 (IRS) |          1.300000e-11|+/-81.E-14  |erg/s/cm^2^         | 8.61E+12|1.300000e+12|                  8.10E+10|                  8.10E+10|                           |                           |+/-8.10E+10    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2010ApJ...709.1257T','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |34.82 microns      |Line measurement; flux integrated over line; lines measured in emission|03 33 36.4 -36 08 25 (J2000)     |Flux integrated from map                                 |LH module                               |From new raw data                                                                                                                                                  
 237|60 microns (IRAS)   |          9.430000e+01|+/-0.033    |Jy                  | 5.00E+12|9.430000e+01|                  3.30E-02|                  3.30E-02|                           |                           |+/-3.30E-02    |Jy       |<a HREF="javascript:getReferenceInfo('2003AJ....126.1607S','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|1 sigma                |60   microns       |Broad-band measurement                                                 |03 33 36.5 -36 08 23 (J2000)     |Total flux                                               |Size, Method, Flag codes: MI;see paper  |From reprocessed raw data                                                                                                                                          
 238|60 microns (ISO)    |          9.200000e+01|+/-20  %    |Jy                  | 5.00E+12|9.200000e+01|                  1.84E+01|                  1.84E+01|                           |                           |+/-1.84E+01    |Jy       |<a HREF="javascript:getReferenceInfo('2001A&A...375..566N','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |60   microns       |Broad-band measurement                                                 |                                 |Modelled datum                                           |                                        |From new raw data                                                                                                                                                  
 241|60 microns (ISO)    |          8.190000e+01|+/-1.0      |Jy                  | 4.93E+12|8.190000e+01|                  1.00E+00|                  1.00E+00|                           |                           |+/-1.00E+00    |Jy       |<a HREF="javascript:getReferenceInfo('2002ApJ...572..105S','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|1 sigma uncert.        |60.8      microns  |Broad-band measurement                                                 |                                 |Flux integrated from map                                 |                                        |From new raw data                                                                                                                                                  
 242|[O I](63) (ISO)     |          5.500000e-15|+/-1.1E-15  |W m^-2^             | 4.76E+12|5.500000e+11|                  1.10E+11|                  1.10E+11|                           |                           |+/-1.10E+11    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2001A&A...375..566N','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |63   microns       |Line measurement; flux integrated over line; lines measured in emission|                                 |Flux integrated from map                                 |                                        |From new raw data                                                                                                                                                  
 243|65 microns (ISO)    |          1.210000e+02|+/-1.0      |Jy                  | 4.45E+12|1.210000e+02|                  1.00E+00|                  1.00E+00|                           |                           |+/-1.00E+00    |Jy       |<a HREF="javascript:getReferenceInfo('2002ApJ...572..105S','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|1 sigma uncert.        |67.3      microns  |Broad-band measurement                                                 |                                 |Flux integrated from map                                 |                                        |From new raw data                                                                                                                                                  
 244|FIR (IRAS)          |          5.070000e-12|            |W m^-2^             | 3.63E+12|1.400000e+02|                          |                          |                           |                           |               |Jy       |<a HREF="javascript:getReferenceInfo('1988ApJS...68...91R','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|82.5 microns       |Broad-band measurement; synthetic band                                 |                                 |Flux integrated from map                                 |                                        |From reprocessed raw data                                                                                                                                          
 245|[O III](88) (ISO)   |          2.700000e-15|+/-0.6E-15  |W m^-2^             | 3.41E+12|2.700000e+11|                  6.00E+10|                  6.00E+10|                           |                           |+/-6.00E+10    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2001A&A...375..566N','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |88   microns       |Line measurement; flux integrated over line; lines measured in emission|                                 |Flux integrated from map                                 |                                        |From new raw data                                                                                                                                                  
 246|90 microns (ISO)    |          1.140000e+02|+/-1.0      |Jy                  | 3.15E+12|1.140000e+02|                  1.00E+00|                  1.00E+00|                           |                           |+/-1.00E+00    |Jy       |<a HREF="javascript:getReferenceInfo('2002ApJ...572..105S','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|1 sigma uncert.        |95.1      microns  |Broad-band measurement                                                 |                                 |Flux integrated from map                                 |                                        |From new raw data                                                                                                                                                  
 247|100 microns (IRAS)  |          1.660000e+02|+/-0.126    |Jy                  | 3.00E+12|1.660000e+02|                  1.26E-01|                  1.26E-01|                           |                           |+/-1.26E-01    |Jy       |<a HREF="javascript:getReferenceInfo('2003AJ....126.1607S','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|1 sigma                |100   microns      |Broad-band measurement                                                 |03 33 36.5 -36 08 23 (J2000)     |Total flux                                               |Size, Method, Flag codes: MI;see paper  |From reprocessed raw data                                                                                                                                          
 250|120 microns (ISO)   |          2.170000e+02|+/-0.80     |Jy                  | 2.52E+12|2.170000e+02|                  8.00E-01|                  8.00E-01|                           |                           |+/-8.00E-01    |Jy       |<a HREF="javascript:getReferenceInfo('2002ApJ...572..105S','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|1 sigma uncert.        |119.0      microns |Broad-band measurement                                                 |                                 |From fitting to map                                      |                                        |From new raw data                                                                                                                                                  
 251|[N II](122) (ISO)   |          2.300000e-15|+/-0.5E-15  |W m^-2^             | 2.46E+12|2.300000e+11|                  5.00E+10|                  5.00E+10|                           |                           |+/-5.00E+10    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2001A&A...375..566N','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |122   microns      |Line measurement; flux integrated over line; lines measured in emission|                                 |Flux integrated from map                                 |                                        |From new raw data                                                                                                                                                  
 252|[C II](158) (ISO)   |          1.100000e-14|+/-2.2E-15  |W m^-2^             | 1.90E+12|1.100000e+12|                  2.20E+11|                  2.20E+11|                           |                           |+/-2.20E+11    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2001A&A...375..566N','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |158   microns      |Line measurement; flux integrated over line; lines measured in emission|                                 |Flux integrated from map                                 |                                        |From new raw data                                                                                                                                                  
 253|150 microns (ISO)   |          1.940000e+02|+/-0.40     |Jy                  | 1.86E+12|1.940000e+02|                  4.00E-01|                  4.00E-01|                           |                           |+/-4.00E-01    |Jy       |<a HREF="javascript:getReferenceInfo('2002ApJ...572..105S','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|1 sigma uncert.        |161.0      microns |Broad-band measurement                                                 |                                 |From fitting to map                                      |                                        |From new raw data                                                                                                                                                  
 254|170 microns (ISO)   |          1.670000e+02|+/-0.60     |Jy                  | 1.72E+12|1.670000e+02|                  6.00E-01|                  6.00E-01|                           |                           |+/-6.00E-01    |Jy       |<a HREF="javascript:getReferenceInfo('2002ApJ...572..105S','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|1 sigma uncert.        |174.0      microns |Broad-band measurement                                                 |                                 |From fitting to map                                      |                                        |From new raw data                                                                                                                                                  
 255|180 microns (ISO)   |          1.030000e+02|+/-0.400    |Jy                  | 1.62E+12|1.030000e+02|                  4.00E-01|                  4.00E-01|                           |                           |+/-4.00E-01    |Jy       |<a HREF="javascript:getReferenceInfo('2002ApJ...572..105S','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|1 sigma uncert.        |185.5      microns |Broad-band measurement                                                 |                                 |From fitting to map                                      |                                        |From new raw data                                                                                                                                                  
 256|200 microns (ISO)   |          8.520000e+01|+/-0.50     |Jy                  | 1.47E+12|8.520000e+01|                  5.00E-01|                  5.00E-01|                           |                           |+/-5.00E-01    |Jy       |<a HREF="javascript:getReferenceInfo('2002ApJ...572..105S','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|1 sigma uncert.        |204.6      microns |Broad-band measurement                                                 |                                 |From fitting to map                                      |                                        |From new raw data                                                                                                                                                  
 257|250 microns (BLAST) |          1.460000e+02|+/-12.9     |Jy                  | 1.20E+12|1.460000e+02|                  1.29E+01|                  1.29E+01|                           |                           |+/-1.29E+01    |Jy       |<a HREF="javascript:getReferenceInfo('2009ApJ...707.1809W','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |250 microns        |Broad-band measurement                                                 |03 33 36.4 -36 08 25 (J2000)     |Total flux                                               |                                        |From new raw data                                                                                                                                                  
 258|350 microns (BLAST) |          6.230000e+01|+/-4.6      |Jy                  | 8.57E+11|6.230000e+01|                  4.60E+00|                  4.60E+00|                           |                           |+/-4.60E+00    |Jy       |<a HREF="javascript:getReferenceInfo('2009ApJ...707.1809W','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |350 microns        |Broad-band measurement                                                 |03 33 36.4 -36 08 25 (J2000)     |Total flux                                               |                                        |From new raw data                                                                                                                                                  
 259|500 microns (BLAST) |          2.470000e+01|+/-2.1      |Jy                  | 6.00E+11|2.470000e+01|                  2.10E+00|                  2.10E+00|                           |                           |+/-2.10E+00    |Jy       |<a HREF="javascript:getReferenceInfo('2009ApJ...707.1809W','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |500 microns        |Broad-band measurement                                                 |03 33 36.4 -36 08 25 (J2000)     |Total flux                                               |                                        |From new raw data                                                                                                                                                  
 261|870 microns (APEX)  |          2.300000e+00|+/-0.3      |Jy                  | 3.45E+11|2.300000e+00|                  3.00E-01|                  3.00E-01|                           |                           |+/-3.00E-01    |Jy       |<a HREF="javascript:getReferenceInfo('2013A&A...555A.128T','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |870 microns        |Broad-band measurement                                                 |03 33 36.37 -36 08 25.4 (J2000)  |Flux integrated from map                                 |                                        |From new raw data                                                                                                                                                  
 262|^12^CO(2-1) (SMA)   |          4.300000e+03|+/-10  %    |Jy km s^-1^         | 2.31E+11|3.290000e+09|                  3.29E+08|                  3.29E+08|                           |                           |+/-3.29E+08    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2007ApJ...654..782S','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |1618   km s^-1^    |Line measurement; flux integrated over line; lines measured in emission|03 33 36.35 -36 08 25.8 (J2000)  |Flux integrated from map                                 |                                        |From new raw data                                                                                                                                                  
 263|^13^CO(2-1) (SMA)   |          3.800000e+02|+/-10  %    |Jy km s^-1^         | 2.20E+11|2.780000e+08|                  2.78E+07|                  2.78E+07|                           |                           |+/-2.78E+07    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2007ApJ...654..782S','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |1618   km s^-1^    |Line measurement; flux integrated over line; lines measured in emission|03 33 36.35 -36 08 25.8 (J2000)  |Flux integrated from map                                 |                                        |From new raw data                                                                                                                                                  
 264|C^18^O(2-1) (SMA)   |          1.100000e+02|+/-10  %    |Jy km s^-1^         | 2.20E+11|8.010000e+07|                  8.01E+06|                  8.01E+06|                           |                           |+/-8.01E+06    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2007ApJ...654..782S','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |1618   km s^-1^    |Line measurement; flux integrated over line; lines measured in emission|03 33 36.35 -36 08 25.8 (J2000)  |Flux integrated from map                                 |                                        |From new raw data                                                                                                                                                  
 265|HC3N 10-9           |                      |<417        |Jy km/s             | 9.10E+10|            |                          |                          |                    1.3E+08|                           |<1.26E+08      |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2011A&A...527A.150L','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|90.979 GHz         |Line measurement; flux integrated over line; lines measured in emission|03 33 36.4 -36 08 26.1 (J2000)   |Flux integrated from map                                 |                                        |From reprocessed raw data                                                                                                                                          
 266|5010 MHz (Parkes)   |          2.100000e-01|+/-0.021    |Jy                  | 5.01E+09|2.100000e-01|                  2.10E-02|                  2.10E-02|                           |                           |+/-2.10E-02    |Jy       |<a HREF="javascript:getReferenceInfo('1970ApL.....5...29W','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|estimated error        |5010       MHz     |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                   |                                        |From new raw data                                                                                                                                                  
 267|5000 MHz            |          1.800000e-01|            |Jy                  | 5.00E+09|1.800000e-01|                          |                          |                           |                           |               |Jy       |<a HREF="javascript:getReferenceInfo('1990PKS90.C...0000W','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|5000   MHz         |Broad-band measurement                                                 |03 31 42.0 -36 18 18 (B1950)     |Integrated from scans                                    |                                        |Homogenized from new and previously published data                                                                                                                 
 268|4.85 GHz (Parkes)   |          2.300000e+02|+/-19       |milliJy             | 4.85E+09|2.300000e-01|                  1.95E-02|                  1.95E-02|                           |                           |+/-1.95E-02    |Jy       |<a HREF="javascript:getReferenceInfo('1996ApJS..103..145W','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|rms noise              |4.85       GHz     |Broad-band measurement                                                 |033340.0 -360824 (J2000)         |Modelled datum                                           |                                        |From new raw data; Corrected for contaminating sources                                                                                                             
 269|4.8 GHz (Effelsberg)|          2.050000e+02|            |milliJy             | 4.80E+09|2.050000e-01|                          |                          |                           |                           |               |Jy       |<a HREF="javascript:getReferenceInfo('2009ApJ...693.1392S','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|4.8 GHz            |Broad-band measurement                                                 |                                 |Flux integrated from map                                 |                                        |From reprocessed raw data                                                                                                                                          
 270|2700 MHz (Parkes)   |          3.400000e-01|            |Jy                  | 2.70E+09|3.400000e-01|                          |                          |                           |                           |               |Jy       |<a HREF="javascript:getReferenceInfo('1990PKS90.C...0000W','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|2700   MHz         |Broad-band measurement                                                 |03 31 42.0 -36 18 18 (B1950)     |Integrated from scans                                    |                                        |Homogenized from new and previously published data                                                                                                                 
 271|1.49 GHz (VLA)      |          5.300000e+02|            |milliJy             | 1.49E+09|5.300000e-01|                          |                          |                           |                           |               |Jy       |<a HREF="javascript:getReferenceInfo('1996ApJS..103...81C','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|1.490   GHz        |Broad-band measurement                                                 |033142.2 -361823 (B1950)         |Total flux                                               |Beamwidth = 48\"                        |Averaged from previously published data                                                                                                                            
 273|HI (21 cm line)     |          1.180000e+01|+/-0.10     |m_21 mag            | 1.42E+09|8.020000e+05|                  7.73E+04|                  7.73E+04|                           |                           |+/-7.73E+04    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('1991RC3.9.C...0000d','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|rms uncertainty        |21         cm      |Line measurement; flux integrated over line; lines measured in emission|033142.0 -361818 (B1950)         |Multiple methods                                         |m_21 equiv. to S(HI) = 8.017E-21 W m^-2 |Homogenized from new and previously published data                                                                                                                 
 274|HI line (Parkes)    |          1.750000e+02|            |Jy km s^-1^         | 1.42E+09|8.230000e+05|                          |                          |                           |                           |               |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2005MNRAS.361...34D','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|1637.1     km s^-1^|Line measurement; flux integrated over line; lines measured in emission|033333.4 -360827. (J2000)        |Flux integrated from map                                 |                                        |Averaged from previously published data                                                                                                                            
 275|HI 21cm line Parkes |          1.460000e+02|+/-8.9      |Jy km/s             | 1.42E+09|6.850000e+05|                  4.18E+04|                  4.18E+04|                           |                           |+/-4.18E+04    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('2004AJ....128...16K','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |1638   km s^-1^    |Line measurement; flux integrated over line                            |03 33 33 -36 08 16 (J2000)       |Flux integrated from map                                 |                                        |From new raw data                                                                                                                                                  
 276|HI (21 cm line)     |          1.350000e+02|+/-10.80    |Jy km s^-1^         | 1.42E+09|6.340000e+05|                  5.07E+04|                  5.07E+04|                           |                           |+/-5.07E+04    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('1989H&RHI.C...0000H','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|21         cm      |Line measurement; flux integrated over line; lines measured in emission|033141.8 -361824. (B1950)        |Not reported in paper                                    |                                        |Transformed from previously published data                                                                                                                         
 277|HI (21 cm line)     |          1.420000e+02|+/-8.00     |Jy km s^-1^         | 1.42E+09|6.670000e+05|                  3.76E+04|                  3.76E+04|                           |                           |+/-3.76E+04    |Jy-Hz    |<a HREF="javascript:getReferenceInfo('1989H&RHI.C...0000H','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|21         cm      |Line measurement; flux integrated over line; lines measured in emission|033141.8 -361824. (B1950)        |Not reported in paper                                    |                                        |Transformed from previously published data                                                                                                                         
 278|HI (21 cm line)     |          1.470000e+02|            |Jy km s^-1^         | 1.42E+09|6.890000e+05|                          |                          |                           |                           |               |Jy-Hz    |<a HREF="javascript:getReferenceInfo('1989H&RHI.C...0000H','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|21         cm      |Line measurement; flux integrated over line; lines measured in emission|033141.8 -361824. (B1950)        |Not reported in paper                                    |                                        |Transformed from previously published data                                                                                                                         
 279|HI (21 cm line)     |          1.960000e+02|            |Jy km s^-1^         | 1.42E+09|9.260000e+05|                          |                          |                           |                           |               |Jy-Hz    |<a HREF="javascript:getReferenceInfo('1996ApJS..107...97M','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|21         cm      |Line measurement; flux integrated over line; lines measured in emission|033141 -361824 (B1950)           |Integrated from scans; Beam filling or dilution corrected|                                        |From new raw data; Corrected for flux in reference beam                                                                                                            
 280|1410 MHz            |          5.300000e-01|            |Jy                  | 1.41E+09|5.300000e-01|                          |                          |                           |                           |               |Jy       |<a HREF="javascript:getReferenceInfo('1990PKS90.C...0000W','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|1410   MHz         |Broad-band measurement                                                 |03 31 42.0 -36 18 18 (B1950)     |Integrated from scans                                    |                                        |Homogenized from new and previously published data                                                                                                                 
 281|1.4GHz              |          3.770000e+02|+/-13.0     |milliJy             | 1.40E+09|3.770000e-01|                  1.30E-02|                  1.30E-02|                           |                           |+/-1.30E-02    |Jy       |<a HREF="javascript:getReferenceInfo('1998AJ....115.1693C','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |1.40   GHz         |Broad-band measurement                                                 |03 33 36.46 -36 08 25.9 (J2000)  |Flux integrated from map                                 |                                        |From new raw data                                                                                                                                                  
 282|843 MHz             |          5.870000e+02|+/-17.7     |milliJy             | 8.43E+08|5.870000e-01|                  1.77E-02|                  1.77E-02|                           |                           |+/-1.77E-02    |Jy       |<a HREF="javascript:getReferenceInfo('2003MNRAS.342.1117M','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |843   MHz          |Broad-band measurement                                                 |033336.41 -360826.1 (J2000)      |Flux integrated from map                                 |                                        |From new raw data                                                                                                                                                  
 283|843 MHz (SUMSS)     |          6.410000e+02|+/-19.3     |milliJy             | 8.43E+08|6.410000e-01|                  1.93E-02|                  1.93E-02|                           |                           |+/-1.93E-02    |Jy       |<a HREF="javascript:getReferenceInfo('2008SUMSS.2.1.....:','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|uncertainty            |843   MHz          |Broad-band measurement                                                 |033336.40 -360826.0 (J2000)      |Flux integrated from map                                 |                                        |From new raw data                                                                                                                                                  
 284|408 MHz (SUMSS)     |          1.060000e+00|+/-0.06     |Jy                  | 4.08E+08|1.060000e+00|                  6.00E-02|                  6.00E-02|                           |                           |+/-6.00E-02    |Jy       |<a HREF="javascript:getReferenceInfo('1981MNRAS.194..693L','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|rms noise              |408        MHz     |Broad-band measurement                                                 |033142.1 -361826 (B1950)         |Modelled datum                                           |                                        |From new raw data; Corrected for contaminating sources                                                                                                             
 285|408 MHz             |          1.060000e+00|            |Jy                  | 4.08E+08|1.060000e+00|                          |                          |                           |                           |               |Jy       |<a HREF="javascript:getReferenceInfo('1990PKS90.C...0000W','_nedInternal');">&nbsp;&nbsp;&nbsp;Ref &swarr;</a>|no uncertainty reported|408   MHz          |Broad-band measurement                                                 |03 31 42.0 -36 18 18 (B1950)     |Integrated from scans                                    |                                        |Homogenized from new and previously published data                                                                                                                 
