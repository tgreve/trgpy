
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-07-07T11:05:25PDT



Photometric Data for GOODS J123702.74+621402.0

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|2-8 keV (Chandra)   ||<-15.85    |log(erg/cm^2^/s)    |1.21E+18||1.17E-11|Jy|2008ApJ...681.1163L|no uncertainty reported|      5.00 keV       | Broad-band measurement|123702.74 +621402.0 (J2000)| Modelled datum|                                        |From reprocessed raw data; NED frequency assigned tomid-point of band in keV
2|0.5-8 keV (Chandra) ||<-16.04    |log(erg/cm^2^/s)    |1.03E+18||8.85E-12|Jy|2008ApJ...681.1163L|no uncertainty reported|      4.25 keV       | Broad-band measurement|123702.74 +621402.0 (J2000)| Modelled datum|                                        |From reprocessed raw data; NED frequency assigned tomid-point of band in keV
3|0.5-2 keV (Chandra) | -16.79    ||log(erg/cm^2^/s)    |3.02E+17|  5.37E-12||Jy|2008ApJ...681.1163L|no uncertainty reported|      1.25 keV       | Broad-band measurement|123702.74 +621402.0 (J2000)| Modelled datum|                                        |From reprocessed raw data; NED frequency assigned tomid-point of band in keV
4|U (KPNO) AB         | 24.6      || mag                |8.22E+14|  5.25E-07||Jy|2004AJ....127.3137C|no uncertainty reported| 3647.65   A         | Broad-band measurement|189.261429 +62.23389 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
5|B F435W (HST/ACS) AB      | 22.558    ||mag                 |6.98E+14|  3.44E-06||Jy|2007ApJ...660...81M|no uncertainty reported|    4297   A         | Broad-band measurement|12 37 02.746 +62 14 01.66 (J2000)| Flux integrated from map|                                        |From reprocessed raw data; Corrected for contaminatingsources
6|B (Subaru) AB       | 24.28     ||mag                 |6.77E+14|  7.05E-07||Jy|2006ApJ...653.1027W|no uncertainty reported| 4427.60   A         | Broad-band measurement|189.261442 62.233794 (J2000)| Flux in fixed aperture|3" diameter aperture                    |Averaged from previously published data
7|B (Subaru) AB       | 24.3      || mag                |6.77E+14|  6.92E-07||Jy|2004AJ....127.3137C|no uncertainty reported| 4427.60   A         | Broad-band measurement|189.261429 +62.23389 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
8|V (Subaru) AB       | 23.9      || mag                |5.48E+14|  1.00E-06||Jy|2004AJ....127.3137C|no uncertainty reported| 5471.22   A         | Broad-band measurement|189.261429 +62.23389 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
9|V (HST/ACS) AB      | 23.094    ||mag                 |5.08E+14|  2.10E-06||Jy|2007ApJ...660...81M|no uncertainty reported|    5907   A         | Broad-band measurement|12 37 02.746 +62 14 01.66 (J2000)| Flux integrated from map|                                        |From reprocessed raw data; Corrected for contaminatingsources
10|R (Keck II) AB      | 23.40     || mag                |4.62E+14|  1.59E-06||Jy|2004AJ....127.3121W|no uncertainty reported|   648.7   A         | Broad-band measurement|12 37 02.746 +62 14 01.66 (J2000)| Total flux|                                        |From new raw data
11|R (Subaru) AB       | 23.20     ||mag                 |4.59E+14|  1.91E-06||Jy|2006ApJ...653.1027W|no uncertainty reported| 6534.16   A         | Broad-band measurement|189.261442 62.233794 (J2000)| Flux in fixed aperture|3" diameter aperture                    |Averaged from previously published data
12|R (Subaru) AB       | 23.2      || mag                |4.59E+14|  1.91E-06||Jy|2004AJ....127.3137C|no uncertainty reported| 6534.16   A         | Broad-band measurement|189.261429 +62.23389 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
13|i F775W (HST/ACS) AB      | 22.499    ||mag                 |3.86E+14|  3.63E-06||Jy|2007ApJ...660...81M|no uncertainty reported|    7764   A         | Broad-band measurement|12 37 02.746 +62 14 01.66 (J2000)| Flux integrated from map|                                        |From reprocessed raw data; Corrected for contaminatingsources
14|I (Subaru) AB       | 22.6      || mag                |3.76E+14|  3.31E-06||Jy|2004AJ....127.3137C|no uncertainty reported| 7975.89   A         | Broad-band measurement|189.261429 +62.23389 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
15|I (Subaru) AB       | 22.62     ||mag                 |3.76E+14|  3.25E-06||Jy|2006ApJ...653.1027W|no uncertainty reported| 7975.89   A         | Broad-band measurement|189.261442 62.233794 (J2000)| Flux in fixed aperture|3" diameter aperture                    |Averaged from previously published data
16|z' (Subaru) AB      | 22.1      || mag                |3.31E+14|  5.25E-06||Jy|2004AJ....127.3137C|no uncertainty reported| 9069.21   A         | Broad-band measurement|189.261429 +62.23389 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
17|z F850LP (HST/ACS) AB      | 21.756    ||mag                 |3.17E+14|  7.21E-06||Jy|2007ApJ...660...81M|no uncertainty reported|    9445   A         | Broad-band measurement|12 37 02.746 +62 14 01.66 (J2000)| Flux integrated from map|                                        |From reprocessed raw data; Corrected for contaminatingsources
18|HK' (QUIRC) AB      | 20.57     |+/-0.05 |mag                 |1.58E+14|  2.15E-05|+/-9.89E-07|Jy|2006ApJ...653.1027W|uncertainty|18947.38   A         | Broad-band measurement|189.261442 62.233794 (J2000)| Flux in fixed aperture|3" diameter aperture                    |Averaged from previously published data
19|HK' (UH) AB         | 20.6      || mag                |1.58E+14|  2.09E-05||Jy|2004AJ....127.3137C|no uncertainty reported|18947.38   A         | Broad-band measurement|189.261429 +62.23389 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
20|3.6 microns (IRAC)  | 55.40     |+/-2.77 |microJy             |8.44E+13|  5.54E-05|+/-2.77E-06|Jy|2011AJ....141....1T|rms uncertainty|     3.550 microns   | Broad-band measurement|189.261414 62.233768 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
21|4.5 microns (IRAC)  | 51.70     |+/-2.59 |microJy             |6.67E+13|  5.17E-05|+/-2.59E-06|Jy|2011AJ....141....1T|rms uncertainty|     4.493 microns   | Broad-band measurement|189.261414 62.233768 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
22|5.8 microns (IRAC)  | 36.70     |+/-1.86 |microJy             |5.23E+13|  3.67E-05|+/-1.86E-06|Jy|2011AJ....141....1T|rms uncertainty|     5.731 microns   | Broad-band measurement|189.261414 62.233768 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
23|8.0 microns (IRAC)  | 44.20     |+/-2.24 |microJy             |3.81E+13|  4.42E-05|+/-2.24E-06|Jy|2011AJ....141....1T|rms uncertainty|     7.872 microns   | Broad-band measurement|189.261414 62.233768 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
24|11 microns (AKARI)  | 61.0      |+/-15   | microJy            |2.73E+13|  6.10E-05|+/-1.50E-05|Jy|2009MNRAS.394..375N|uncertainty|        11 microns   | Broad-band measurement|12 37 02.74 +62 14 02.02 (J2000)| Flux integrated from map|                                        |From new raw data
25|ISOCAM 15 microns   | 0.3322    |+/-0.1  |milliJy             |2.07E+13|  3.32E-04|+/-1.00E-04|Jy|1997MNRAS.289..465G|estimated error|14.5       microns   | Broad-band measurement|123702.57 +621406.1 (J2000)| Flux integrated from map|                                        |From new raw data
26|15 microns (ISOCAM) | 144       |+/-20   |microJy             |2.00E+13|  1.44E-04|+/-2.00E-05|Jy|2006A&A...451...57M|68% confidence|    15.0   microns   | Broad-band measurement|189.2614288 62.2338943 (J2000)| Flux integrated from map|                                        |Averaged from previously published data
27|16 microns (IRS)    | 441.9     |+/-17.8 |microJy             |1.90E+13|  4.42E-04|+/-1.78E-05|Jy|2011AJ....141....1T|rms uncertainty|      15.8 microns   | Broad-band measurement|189.261414 62.233768 (J2000)| From fitting to map|                                        |From new raw data
28|18 microns (AKARI)  | 417       |+/-33   | microJy            |1.67E+13|  4.17E-04|+/-3.30E-05|Jy|2009MNRAS.394..375N|uncertainty|        18 microns   | Broad-band measurement|12 37 02.74 +62 14 02.02 (J2000)| Flux integrated from map|                                        |From new raw data
29|24 microns (MIPS)   | 349.0     |+/-8.8  |microJy             |1.27E+13|  3.49E-04|+/-8.80E-06|Jy|2011AJ....141....1T|rms uncertainty|     23.68 microns   | Broad-band measurement|189.261414 62.233768 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
30|24 microns (MIPS)   | 347.3     |+/-4.5  |microJy             |1.27E+13|  3.47E-04|+/-4.50E-06|Jy|2011A&A...528A..35M|uncertainty|     23.68 microns   | Broad-band measurement|12 37 02.74 +62 14 01.50 (J2000)| Flux integrated from map|                                        |From new raw data
31|24 microns (MIPS)   | 334       |+/-8    |microJy             |1.27E+13|  3.34E-04|+/-8.00E-06|Jy|2006A&A...451...57M|68% confidence|   23.68   microns   | Broad-band measurement|189.2614288 62.2338943 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
32|70 microns (MIPS)   | 2.6       |+/-0.2  |milliJy             |4.20E+12|  2.60E-03|+/-2.00E-04|Jy|2011A&A...528A..35M|uncertainty|     71.42 microns   | Broad-band measurement|12 37 02.74 +62 14 01.50 (J2000)| Flux integrated from map|                                        |From new raw data
33|1.4 GHz (VLA)       | 40        |+/-12   | microJy            |1.40E+09|  4.00E-05|+/-1.20E-05|Jy|2006MNRAS.371..963B|1 sigma|       1.4 GHz       | Broad-band measurement|12 37 02.710 +62 14 01.84 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
34|1.4 GHz (VLA)       | 41.1      |+/-7.8  |microJy             |1.40E+09|  4.11E-05|+/-7.80E-06|Jy|2010ApJS..188..178M|uncertainty|       1.4 GHz       | Broad-band measurement|12 37 02.73 +62 14 01.6 (J2000)| Total flux; Beam filling or dilution corrected|Major=1.1"; Minor=0.0"; PA=121 deg      |From new raw data
35|1.4 GHz (VLA)       | 30.39     ||microJy             |1.40E+09|  3.04E-05||Jy|2006A&A...451...57M|no uncertainty reported|     1.4   GHz       | Broad-band measurement|189.2614288 62.2338943 (J2000)| Flux integrated from map|                                        |From new raw data
