
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-07-10T13:09:38PDT



Photometric Data for B2 2327+39

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|3.6 microns (IRAC)  | 99.6      |+/-10.1 | microJy            |8.44E+13|  9.96E-05|+/-1.01E-05|Jy|2007ApJS..171..353S|uncertainty|   3.550   microns   | Broad-band measurement|23 30 24.9 +39 27 12.02 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
2|4.5 microns (IRAC)  | 143.0     |+/-14.0 | microJy            |6.67E+13|  1.43E-04|+/-1.40E-05|Jy|2007ApJS..171..353S|uncertainty|   4.493   microns   | Broad-band measurement|23 30 24.9 +39 27 12.02 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
3|5.8 microns (IRAC)  | 160.0     |+/-16.0 | microJy            |5.23E+13|  1.60E-04|+/-1.60E-05|Jy|2007ApJS..171..353S|uncertainty|   5.731   microns   | Broad-band measurement|23 30 24.9 +39 27 12.02 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
4|8.0 microns (IRAC)  | 474.0     |+/-47.0 | microJy            |3.81E+13|  4.74E-04|+/-4.70E-05|Jy|2007ApJS..171..353S|uncertainty|   7.872   microns   | Broad-band measurement|23 30 24.9 +39 27 12.02 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
5|16 microns (IRS)    | 1040.0    |+/-88.0 | microJy            |1.87E+13|  1.04E-03|+/-8.80E-05|Jy|2007ApJS..171..353S|uncertainty|      16   microns   | Broad-band measurement|23 30 24.9 +39 27 12.02 (J2000)| Flux in fixed aperture|6" diameter aperture                    |From reprocessed raw data
6|24 microns (MIPS)   | 2210.0    |+/-113.2| microJy            |1.27E+13|  2.21E-03|+/-1.13E-04|Jy|2007ApJS..171..353S|uncertainty|   23.68   microns   | Broad-band measurement|23 30 24.9 +39 27 12.02 (J2000)| Flux in fixed aperture|13" diameter aperture                   |From reprocessed raw data
7|70 microns (MIPS)   ||<4670      | microJy            |4.20E+12||4.67E-03|Jy|2007ApJS..171..353S|3 sigma|   71.42   microns   | Broad-band measurement|23 30 24.9 +39 27 12.02 (J2000)| Flux in fixed aperture|35" diameter aperture                   |From reprocessed raw data
3|100 microns (PACS) | 11.3       |+/-2.9  |mJy             |2.998e+12| 11.3E-03 |+/-2.9E-03|Jy|2005MNRAS.358..149P|1rms uncertainty|     850   microns   | Broad-band measurement|12 37 11.7 +62 22 12 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
4|160 microns (PACS) | 27.0     |+/-6.2 |mJy             |1.874e+12| 27.0E-03|+/-6.2E-03 |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
8|160 microns (MIPS)  ||<64300     | microJy            |1.92E+12||6.43E-02|Jy|2007ApJS..171..353S|3 sigma|   155.9   microns   | Broad-band measurement|23 30 24.9 +39 27 12.02 (J2000)| Flux in fixed aperture|50" diameter aperture                   |From reprocessed raw data
5|250 microns (SPIRE)| 52.      |+/-2.7 |mJy             |1.199e+12| 52.0E-03|+/-2.7e-03 |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
6|350 microns (SPIRE)| 60.3      |+/-2.7  |mJy             |8.565e+11|60.3E-03 |+/-2.7e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
8|500 microns (SPIRE) | 57.3     |+/-3.3 |mJy             |5.996e+11|57.3E-03 |+/-3.3e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
9|450 microns (SCUBA) | 49        |+/-18   | milliJy            |6.66E+11|  4.90E-02|+/-1.80E-02|Jy|2004MNRAS.353..377R|uncertainty|       450 microns   | Broad-band measurement|23 30 24.91 +39 27 11.2 (J2000)| Not reported in paper|Good quality data                       |From new raw data
10|850 microns (SCUBA) | 14.1      |+/-1.7  | milliJy            |3.53E+11|  1.41E-02|+/-1.70E-03|Jy|2004MNRAS.353..377R|uncertainty|       850 microns   | Broad-band measurement|23 30 24.91 +39 27 11.2 (J2000)| Not reported in paper|Good quality data                       |From new raw data
10|850 microns (SCUBA) | 22.2      |+/-2.7  | milliJy            |3.53E+11|  22.2E-03|+/-2.7E-03|Jy|2004MNRAS.353..377R|uncertainty|       850 microns   | Broad-band measurement|23 30 24.91 +39 27 11.2 (J2000)| Not reported in paper|Good quality data                       |From new raw data
11|4.85 GHz            | 34        |+/-6    |milliJy             |4.85E+09|  3.40E-02|+/-6.00E-03|Jy|1991ApJS...75.1011G|rms noise|4.85       GHz       | Broad-band measurement|232800.5 +391033 (B1950)| Modelled datum|                                        |From new raw data; Corrected for contaminating sources
12|4.85 GHz            | 32        |+/-15  %|milliJy             |4.85E+09|  3.20E-02|+/-4.80E-03|Jy|1991ApJS...75....1B|uncertainty|4.85       GHz       | Broad-band measurement|232800.6 +391041 (B1950)| Peak flux|                                        |From new raw data; Corrected for contaminating sources
13|1.4GHz (VLA)        | 100.0     |+/-3.0  |milliJy             |1.40E+09|  1.00E-01|+/-3.00E-03|Jy|1998AJ....115.1693C|uncertainty|    1.40   GHz       | Broad-band measurement|23 30 24.91 +39 27 11.5 (J2000)| Flux integrated from map|                                        |From new raw data
14|408 MHz             | 0.36      |+/-0.02 |Jy                  |4.08E+08|  3.60E-01|+/-2.13E-02|Jy|1985A&AS...59..255F|rms uncertainty|408        MHz       | Broad-band measurement|23 27 59.7 39 10 54 (B1950)| Total flux|                                        |From new raw data
15|408 MHz             | 0.269     |+/-0.07 |Jy                  |4.08E+08|  2.69E-01|+/-7.00E-02|Jy|1973A&AS...11..291C|internal error|408        MHz       | Broad-band measurement; peak value reported|232757.8 +390954. (B1950)| Peak flux|                                        |From new raw data
16|365 MHz (Texas)     | 0.394     |+/-0.023|Jy                  |3.65E+08|  3.94E-01|+/-2.30E-02|Jy|1996AJ....111.1945D|internal error|365        MHz       | Broad-band measurement; obtained by interpolation over frequency|232758.404 391038.98 (B1950)| Integrated from scans|Model:P;MFlag:+;EFlag:+;LFlag:C.        |From new raw data
17|74 MHz (VLA)        | 1.74      |+/-0.20 | Jy                 |7.38E+07|  1.74E+00|+/-2.00E-01|Jy|2007AJ....134.1245C|rms uncertainty|      73.8 MHz       | Broad-band measurement|23 30 25.09 +39 27 09.3 (J2000)| Flux integrated from map|Corrected for clean bias                |From new raw data
