
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-12-12T09:48:50PST



Photometric Data for SMM J041327.2+102743

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|3.6 microns (IRAC)  | 6.2415E+01|+/-3.9744E-01|microJy             |8.44E+13|  6.24E-05|+/-3.97E-07|Jy|2013SSTSLC4.2....0C|uncertainty|3.55       microns   | Broad-band measurement|| Flux in fixed aperture|5.8" aperture                           |From new raw data
2|3.6 microns (IRAC)  | 5.6688E+01|+/-2.7508E-01|microJy             |8.44E+13|  5.67E-05|+/-2.75E-07|Jy|2013SSTSLC4.2....0C|uncertainty|3.55       microns   | Broad-band measurement|| Flux in fixed aperture|3.8" aperture                           |From new raw data
3|4.5 microns (IRAC)  | 8.6521E+01|+/-4.0974E-01|microJy             |6.67E+13|  8.65E-05|+/-4.10E-07|Jy|2013SSTSLC4.2....0C|uncertainty|4.493      microns   | Broad-band measurement|| Flux in fixed aperture|3.8" aperture                           |From new raw data
4|4.5 microns (IRAC)  | 9.2896E+01|+/-6.0378E-01|microJy             |6.67E+13|  9.29E-05|+/-6.04E-07|Jy|2013SSTSLC4.2....0C|uncertainty|4.493      microns   | Broad-band measurement|| Flux in fixed aperture|5.8" aperture                           |From new raw data
5|5.8 microns (IRAC)  | 1.4492E+02|+/-1.7675E+00|microJy             |5.23E+13|  1.45E-04|+/-1.77E-06|Jy|2013SSTSLC4.2....0C|uncertainty|5.731      microns   | Broad-band measurement|| Flux in fixed aperture|3.8" aperture                           |From new raw data
6|5.8 microns (IRAC)  | 1.4808E+02|+/-2.4772E+00|microJy             |5.23E+13|  1.48E-04|+/-2.48E-06|Jy|2013SSTSLC4.2....0C|uncertainty|5.731      microns   | Broad-band measurement|| Flux in fixed aperture|5.8" aperture                           |From new raw data
7|8.0 microns (IRAC)  | 3.5606E+02|+/-3.7470E+00|microJy             |3.81E+13|  3.56E-04|+/-3.75E-06|Jy|2013SSTSLC4.2....0C|uncertainty|7.872      microns   | Broad-band measurement|| Flux in fixed aperture|5.8" aperture                           |From new raw data
8|8.0 microns (IRAC)  | 3.6087E+02|+/-2.8295E+00|microJy             |3.81E+13|  3.61E-04|+/-2.83E-06|Jy|2013SSTSLC4.2....0C|uncertainty|7.872      microns   | Broad-band measurement|| Flux in fixed aperture|3.8" aperture                           |From new raw data
9|24 microns (MIPS)   | 1.4939E+03|+/-3.4580E+01|microJy             |1.27E+13|  1.49E-03|+/-3.46E-05|Jy|2013SSTSLC4.2....0C|uncertainty|23.68      microns   | Broad-band measurement|| Modelled datum|PSF fit                                 |From new raw data
10|24 microns (MIPS)   | 1.5003E+03|+/-3.1890E+01|microJy             |1.27E+13|  1.50E-03|+/-3.19E-05|Jy|2013SSTSLC4.2....0C|uncertainty|23.68      microns   | Broad-band measurement|| Flux in fixed aperture|14.7" aperture                          |From new raw data
11|450 microns (SCUBA) | 55.4      |+/-16.6 | milliJy            |6.66E+11|  5.54E-02|+/-1.66E-02|Jy|2008MNRAS.384.1611K|rms uncertainty|       450 microns   | Broad-band measurement|041327.2 +102743 (J2000)| Flux integrated from map|S/N = 5.3                               |From new raw data
12|450 microns (SCUBA) | 11        |+/-33   |milliJy             |6.66E+11|  1.10E-02|+/-3.30E-02|Jy|2007MNRAS.376.1073Z|uncertainty|     450   microns   | Broad-band measurement|04 13 26.9 +10 27 41 (J2000)| Flux integrated from map|                                        |From reprocessed raw data
13|850 microns (SCUBA) | 30.0      ||milliJy             |3.53E+11|  3.00E-02||Jy|2007MNRAS.376.1073Z|no uncertainty reported|     850   microns   | Broad-band measurement|04 13 26.9 +10 27 41 (J2000)| Flux integrated from map|S/N = 16.2                              |From reprocessed raw data
14|850 microns (SCUBA) | 25.0      |+/-2.8  | milliJy            |3.53E+11|  2.50E-02|+/-2.80E-03|Jy|2008MNRAS.384.1611K|rms uncertainty|       850 microns   | Broad-band measurement|041327.2 +102743 (J2000)| Flux integrated from map|S/N = 14.4                              |From new raw data
14|3mm OVRO            |           |<0.9  | milliJy            |99.9E+9|  |0.9E-03|Jy|2008MNRAS.384.1611K|3sigma uncertainty|       850 microns   | Broad-band measurement|041327.2 +102743 (J2000)| Flux integrated from map|S/N = 14.4                              |From new raw data
15|CO(3-2) (OVRO)      | 5.4       |+/-1.3  | Jy km/s            |3.46E+11|  1.62E+06|+/-3.90E+05|Jy-Hz|2004ApJ...609...61H|uncertainty|   2.846             | Line measurement; flux integrated over line; lines measured in emission|04 13 27.50 +10 27 40.3 (J2000)| Flux integrated from map|                                        |From new raw data
16|CO(1-0) (GBT)       | 0.644     |+/-0.082|Jy km/s             |1.15E+11|  6.44E+04|+/-8.19E+03|Jy-Hz|2011ApJ...739L..32R|uncertainty|   115.271 GHz       | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|Measured with Spectrometer backend      |From new raw data
14|1.4 GHz (VLA)       |           |<1.5| milliJy            |1.40E+11| |1.5E-03|Jy|2004A&A...423..441B|3sigma uncertainty|    1.4    GHz       | Broad-band measurement|14 09 55.57 +56 28 26.47 (J2000)| Flux integrated from map|                                        |From new raw data
