
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-06-16T17:15:19PDT



Photometric Data for [HB89] 2343+125:MD0059

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|G (WHT)             | 24.99     ||mag                 |6.38E+14|  3.67E-07||Jy|2006ApJ...647..128E|no uncertainty reported|    0.47   microns   | Broad-band measurement|| Flux in fixed aperture|                                        |Averaged from previously published data
2|R (Hale)            | 24.99     || mag                |4.76E+14|  3.11E-07||Jy|2007ApJ...670...15R|no uncertainty reported|      6300 A         | Broad-band measurement|| Not reported in paper|                                        |Averaged new and previously published data
3|H{alpha} (Keck II)  | 2.9E-17   |+/-0.4E-17|erg s^-1^ cm^-2^    |4.57E+14|  2.90E+06|+/-4.00E+05|Jy-Hz|2006ApJ...646..107E|uncertainty|    6563   A         | Line measurement; flux integrated over line; lines measured in emission|23 46 26.90 +12 47 39.87 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
4|J (Hale/WIRC)       | 22.73     ||mag                 |2.40E+14|  1.26E-06||Jy|2006ApJ...646..107E|no uncertainty reported|    1.25   microns   | Broad-band measurement|23 46 26.90 +12 47 39.87 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data; derived from aflux in a different band and a color
5|K_s (Hale/WIRC)     | 20.14     ||mag                 |1.39E+14|  5.89E-06||Jy|2006ApJ...646..107E|no uncertainty reported|    2.15   microns   | Broad-band measurement|23 46 26.90 +12 47 39.87 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data
