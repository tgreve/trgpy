
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-07-10T13:42:15PDT



Photometric Data for SPT-S J045912-5942.4

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|1.4 mm (SPT)        | 20.85     |+/-3.90 |milliJy             |2.20E+11|  2.09E-02|+/-3.90E-03|Jy|2010ApJ...719..763V|uncertainty|       1.4 mm        | Broad-band measurement|74.804 -59.708 (J2000)| Flux integrated from map|De-boosted flux; S/N = 7.05             |From new raw data
2|1.4 mm (SPT)        | 22.58     ||milliJy             |2.20E+11|  2.26E-02||Jy|2010ApJ...719..763V|no uncertainty reported|       1.4 mm        | Broad-band measurement|74.804 -59.708 (J2000)| Flux integrated from map|Raw flux; S/N = 7.05                    |From new raw data
3|2.0 mm (SPT)        | 7.26      |+/-1.27 |milliJy             |1.50E+11|  7.26E-03|+/-1.27E-03|Jy|2010ApJ...719..763V|uncertainty|       2.0 mm        | Broad-band measurement|74.804 -59.708 (J2000)| Flux integrated from map|De-boosted flux; S/N = 6.20             |From new raw data
4|2.0 mm (SPT)        | 7.51      ||milliJy             |1.50E+11|  7.51E-03||Jy|2010ApJ...719..763V|no uncertainty reported|       2.0 mm        | Broad-band measurement|74.804 -59.708 (J2000)| Flux integrated from map|Raw flux; S/N = 6.20                    |From new raw data
