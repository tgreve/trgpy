
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-04-05T06:04:16PDT



Photometric Data for SMM J163555.5+661300

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|450 microns (SCUBA) | 18.0      |+/-5.4  |milliJy             |6.66E+11|  1.80E-02|+/-5.40E-03|Jy|2006MNRAS.368..487K|uncertainty|     450   microns   | Broad-band measurement|163555.5 +661300 (J2000)| Flux integrated from map|                                        |From new raw data
2|450 microns (SCUBA) | 2         |+/-25   |milliJy             |6.66E+11|  2.00E-03|+/-2.50E-02|Jy|2007MNRAS.376.1073Z|uncertainty|     450   microns   | Broad-band measurement|16 35 55.5 +66 12 58 (J2000)| Flux integrated from map|                                        |From reprocessed raw data
3|450 microns (SCUBA) | |<11.8      | milliJy            |6.66E+11| |1.18E-02|Jy|2008MNRAS.384.1611K|1sigma uncertainty reported|       450 microns   | Broad-band measurement|163555.5 +661300 (J2000)| Flux integrated from map|                                        |From new raw data
4|CO(4-3) (IRAM)      | |<0.45      | Jy km/s            |4.61E+11| |5.89E-08|Jy|2009A&A...496...45K|3 sigma|   461.041 GHz       | Line measurement; flux integrated over line; lines measured in emission|16 35 56.01 +66 12 54.3 (J2000)| Flux integrated from map|                                        |From new raw data
5|850 microns (SCUBA) | 11.3      |+/-1.3  | milliJy            |3.53E+11|  1.13E-02|+/-1.30E-03|Jy|2008MNRAS.384.1611K|rms uncertainty|       850 microns   | Broad-band measurement|163555.5 +661300 (J2000)| Flux integrated from map|S/N = 15.8                              |From new raw data
6|850 microns (SCUBA) | 6.2       | |milliJy             |3.53E+11|  6.20E-03| |Jy|2007MNRAS.376.1073Z|no uncertainty reported|     850   microns   | Broad-band measurement|16 35 55.5 +66 12 58 (J2000)| Flux integrated from map|S/N = 8.7                               |From reprocessed raw data
7|850 microns (SCUBA) | 11.3      |+/-1.3  |milliJy             |3.53E+11|  1.13E-02|+/-1.30E-03|Jy|2006MNRAS.368..487K|uncertainty|     850   microns   | Broad-band measurement|163555.5 +661300 (J2000)| Flux integrated from map|                                        |From new raw data
8|870 microns (SMA)   | 10.7      |+/-2.0  |milliJy             |3.40E+11|  1.07E-02|+/-2.00E-03|Jy|2010ApJ...709..210K|uncertainty|      870  microns   | Broad-band measurement|16 35 55.67 +66 12 59.51 (J2000)| Flux integrated from map|                                        |From new raw data
9|3 mm (IRAM)         | |<0.44      | milliJy            |9.99E+10| |4.40E-04|Jy|2009A&A...496...45K|3sigma uncertainty|         3 mm        | Broad-band measurement|16 35 56.01 +66 12 54.3 (J2000)| Flux integrated from map|                                        |From new raw data
