
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-05-30T03:36:06PDT



Photometric Data for RG J131208.34+424144.4

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|R (SUBARU)          | 23.4      |+/-0.3  |mag                 |4.76E+14|  1.36E-06|+/-3.76E-07|Jy|2006ApJS..167..103F|rms uncertainty|    6300   A         | Broad-band measurement|| Flux in fixed aperture|3" radius aperture                      |From new raw data
4|I (Cousins)         | 22.91     |+/-0.04 |mag                 |3.79E+14|  1.75E-06|+/-6.56E-08|Jy|2004ApJ...616...71S|1 sigma|    7900   A         | Broad-band measurement|| Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
5|z (SUBARU)          | 22.4      |+/-0.5  |mag                 |3.26E+14|  2.40E-06|+/-1.11E-06|Jy|2006ApJS..167..103F|rms uncertainty|    9200   A         | Broad-band measurement|| Flux in fixed aperture|3" radius aperture                      |From new raw data
6|J (2MASS)           | 22.92     |+/-0.30 |mag                 |2.40E+14|  1.08E-06|+/-3.44E-07|Jy|2004ApJ...616...71S|1 sigma|    1.25   microns   | Broad-band measurement|| Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
7|K_s_ (2MASS)        | 19.10     |+/-0.12 |mag                 |1.38E+14|  1.53E-05|+/-1.79E-06|Jy|2004ApJ...616...71S|1 sigma|    2.17   microns   | Broad-band measurement|| Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
1|24 microns (MIPS)   | 279       |+/-14   |mJy                 |1.27E+13|279.E-06|14.0E-06|Jy|2009ApJ...694.1517D|3sigma uncertainty|     23.68 microns   | Broad-band measurement|12 37 11.89 +62 22 11.8 (J2000)| Flux integrated from map|                                        |From new raw data
2|350 microns (SPIRE) |           |<82     |mJy                 |8.565e+11||82.0e-03       |Jy|2.40e+01           |3sigma uncertainty|-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
8|850 microns (SCUBA) | 1.8       |+/-1.5  | milliJy            |3.53E+11|  1.80E-03|+/-1.50E-03|Jy|2004ApJ...614..671C|uncertainty|       850 microns   | Broad-band measurement|131208.34 +424144.4 (J2000)| Flux integrated from map|                                        |From new raw data
8|850 microns (SCUBA) |        |<4.5  | milliJy            |3.53E+11|  |4.5E-03|Jy|2004ApJ...614..671C|3sigma uncertainty|       850 microns   | Broad-band measurement|131208.34 +424144.4 (J2000)| Flux integrated from map|                                        |From new raw data
9|1.4 GHz (VLA)       | 37        |+/-15   |microJy             |1.40E+09|  3.70E-05|+/-1.50E-05|Jy|2006ApJS..167..103F|uncertainty|     1.4   GHz       | Broad-band measurement|13 12 08.367 +42 41 44.77 (J2000)| Flux integrated from map|Corrected to the sky; see paper         |From new raw data
9|1.4 GHz (VLA)       | 37.6        |+/-4.0   |microJy             |1.40E+09|  3.76E-05|+/-4.00E-06|Jy|2006ApJS..167..103F|uncertainty|     1.4   GHz       | Broad-band measurement|13 12 08.367 +42 41 44.77 (J2000)| Flux integrated from map|Corrected to the sky; see paper         |From new raw data
