
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-07-10T07:03:41PDT



Photometric Data for BRI 1335-0417

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
2|350 microns (SHARC-II)        | 0.052     |+/-0.008|Jy                  |8.57E+11|  5.20E-02|+/-8.00E-03|Jy|1999CIT...T00R....B|1 sigma|350        microns   | Broad-band measurement|133527.6 -041721. (B1950)| Flux integrated from map|                                        |From new raw data
5|1.4 GHz (VLBI)      | 208       |+/-46   | microJy            |1.40E+09|  2.08E-04|+/-4.60E-05|Jy|2007AJ....134..694M|uncertainty|    1.4    GHz       | Broad-band measurement|| Total flux|                                        |From new raw data
