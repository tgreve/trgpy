
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-07-10T07:33:59PDT



Photometric Data for 2MASSi J1649149+530316

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|H{alpha} (TNG)      | 3.1E-14   |+/-20  %|erg/s/cm^2^         |4.57E+14|  3.10E+09|+/-6.20E+08|Jy-Hz|2011A&A...531A.128O|uncertainty|      6563 A         | Line measurement; flux integrated over line; lines measured in emission|16 49 14 +53 03 16 (J2000)| From fitting to map|Broad component flux                    |From new raw data
2|H{alpha} (TNG)      | 2.3E-14   |+/-20  %|erg/s/cm^2^         |4.57E+14|  2.30E+09|+/-4.60E+08|Jy-Hz|2011A&A...531A.128O|uncertainty|      6563 A         | Line measurement; flux integrated over line; lines measured in emission|16 49 14 +53 03 16 (J2000)| From fitting to map|Intermediate component flux             |From new raw data
3|6.7 microns (IRS)   | 9.4       || milliJy            |4.47E+13|  9.40E-03||Jy|2007A&A...468..979M|no uncertainty reported|     6.7   microns   | Broad-band measurement|16 49 14.90 +53 03 16.0 (J2000)| Flux integrated from map|                                        |From new raw data
4|250 GHz (IRAM/MAMBO)| 4.6E-03   |+/-0.8E-03|Jy                  |2.50E+11|  4.60E-03|+/-8.00E-04|Jy|2006AJ....132.1307P|1 sigma|     250   GHz       | Broad-band measurement|16 49 15.02 +53 03 16.5 (J2000)| Flux integrated from map|From 2003A&A...398..857O                |Averaged from previously published data
5|5.0 GHz (VLA)       | 910E-06   |+/-80E-06|Jy                  |5.00E+09|  9.10E-04|+/-8.00E-05|Jy|2006AJ....132.1307P|1 sigma|     5.0   GHz       | Broad-band measurement|16 49 15.02 +53 03 16.5 (J2000)| Flux integrated from map|                                        |From new raw data
6|1.4 GHz (VLA)       | 820E-06   |+/-20E-06|Jy                  |1.40E+09|  8.20E-04|+/-2.00E-05|Jy|2006AJ....132.1307P|1 sigma|     1.4   GHz       | Broad-band measurement|16 49 15.02 +53 03 16.5 (J2000)| Flux integrated from map|                                        |From new raw data
