
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-07-08T04:27:48PDT



Photometric Data for GOODS J123709.14+621508.3

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|B F435W (HST/ACS) AB      | 23.805    ||mag                 |6.98E+14|  1.09E-06||Jy|2007ApJ...660...81M|no uncertainty reported|    4297   A         | Broad-band measurement|12 37 09.128 +62 15 07.91 (J2000)| Flux integrated from map|                                        |From reprocessed raw data; Corrected for contaminatingsources
2|B (Subaru) AB       | 23.95     ||mag                 |6.77E+14|  9.55E-07||Jy|2006ApJ...653.1027W|no uncertainty reported| 4427.60   A         | Broad-band measurement|189.288033 62.252197 (J2000)| Flux in fixed aperture|3" diameter aperture                    |Averaged from previously published data
3|V (HST/ACS) AB      | 23.399    ||mag                 |5.08E+14|  1.59E-06||Jy|2007ApJ...660...81M|no uncertainty reported|    5907   A         | Broad-band measurement|12 37 09.128 +62 15 07.91 (J2000)| Flux integrated from map|                                        |From reprocessed raw data; Corrected for contaminatingsources
4|R (Keck II) AB      | 23.51     || mag                |4.62E+14|  1.43E-06||Jy|2004AJ....127.3121W|no uncertainty reported|   648.7   A         | Broad-band measurement|12 37 09.128 +62 15 07.91 (J2000)| Total flux|                                        |From new raw data
5|R (Subaru) AB       | 23.25     ||mag                 |4.59E+14|  1.82E-06||Jy|2006ApJ...653.1027W|no uncertainty reported| 6534.16   A         | Broad-band measurement|189.288033 62.252197 (J2000)| Flux in fixed aperture|3" diameter aperture                    |Averaged from previously published data
6|i F775W (HST/ACS) AB      | 22.759    ||mag                 |3.86E+14|  2.86E-06||Jy|2007ApJ...660...81M|no uncertainty reported|    7764   A         | Broad-band measurement|12 37 09.128 +62 15 07.91 (J2000)| Flux integrated from map|                                        |From reprocessed raw data; Corrected for contaminatingsources
7|I (Subaru) AB       | 22.75     ||mag                 |3.76E+14|  2.88E-06||Jy|2006ApJ...653.1027W|no uncertainty reported| 7975.89   A         | Broad-band measurement|189.288033 62.252197 (J2000)| Flux in fixed aperture|3" diameter aperture                    |Averaged from previously published data
8|z F850LP (HST/ACS) AB      | 22.069    ||mag                 |3.17E+14|  5.40E-06||Jy|2007ApJ...660...81M|no uncertainty reported|    9445   A         | Broad-band measurement|12 37 09.128 +62 15 07.91 (J2000)| Flux integrated from map|                                        |From reprocessed raw data; Corrected for contaminatingsources
9|HK' (QUIRC) AB      | 21.04     |+/-0.12 |mag                 |1.58E+14|  1.39E-05|+/-1.54E-06|Jy|2006ApJ...653.1027W|uncertainty|18947.38   A         | Broad-band measurement|189.288033 62.252197 (J2000)| Flux in fixed aperture|3" diameter aperture                    |Averaged from previously published data
10|3.6 microns (IRAC)  | 26.40     |+/-0.04 |microJy             |8.44E+13|  2.64E-05|+/-4.00E-08|Jy|2009ApJ...705...68B|uncertainty|     3.550 microns   | Broad-band measurement|189.288 62.2524 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
11|3.6 microns (IRAC)  | 27.00     |+/-1.35 |microJy             |8.44E+13|  2.70E-05|+/-1.35E-06|Jy|2011AJ....141....1T|rms uncertainty|     3.550 microns   | Broad-band measurement|189.288086 62.252220 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
12|4.5 microns (IRAC)  | 24.50     |+/-0.06 |microJy             |6.67E+13|  2.45E-05|+/-6.00E-08|Jy|2009ApJ...705...68B|uncertainty|     4.493 microns   | Broad-band measurement|189.288 62.2524 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
13|4.5 microns (IRAC)  | 24.90     |+/-1.25 |microJy             |6.67E+13|  2.49E-05|+/-1.25E-06|Jy|2011AJ....141....1T|rms uncertainty|     4.493 microns   | Broad-band measurement|189.288086 62.252220 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
14|5.8 microns (IRAC)  | 18.50     |+/-0.32 |microJy             |5.23E+13|  1.85E-05|+/-3.20E-07|Jy|2009ApJ...705...68B|uncertainty|     5.731 microns   | Broad-band measurement|189.288 62.2524 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
15|5.8 microns (IRAC)  | 18.20     |+/-0.97 |microJy             |5.23E+13|  1.82E-05|+/-9.70E-07|Jy|2011AJ....141....1T|rms uncertainty|     5.731 microns   | Broad-band measurement|189.288086 62.252220 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
16|8.0 microns (IRAC)  | 17.90     |+/-0.35 |microJy             |3.81E+13|  1.79E-05|+/-3.50E-07|Jy|2009ApJ...705...68B|uncertainty|     7.872 microns   | Broad-band measurement|189.288 62.2524 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
17|8.0 microns (IRAC)  | 18.10     |+/-0.99 |microJy             |3.81E+13|  1.81E-05|+/-9.90E-07|Jy|2011AJ....141....1T|rms uncertainty|     7.872 microns   | Broad-band measurement|189.288086 62.252220 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
18|16 microns (IRS)    | 142.0     |+/-7.8  |microJy             |1.90E+13|  1.42E-04|+/-7.80E-06|Jy|2011AJ....141....1T|rms uncertainty|      15.8 microns   | Broad-band measurement|189.288086 62.252220 (J2000)| From fitting to map|                                        |From new raw data
19|24 microns (MIPS)   | 123.0     |+/-5.4  |microJy             |1.27E+13|  1.23E-04|+/-5.40E-06|Jy|2009ApJ...705...68B|uncertainty|     23.68 microns   | Broad-band measurement|189.288 62.2524 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
20|24 microns (MIPS)   | 123.0     |+/-5.8  |microJy             |1.27E+13|  1.23E-04|+/-5.80E-06|Jy|2011AJ....141....1T|rms uncertainty|     23.68 microns   | Broad-band measurement|189.288086 62.252220 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
21|24 microns (MIPS)   | 127.8     |+/-2.7  |microJy             |1.27E+13|  1.28E-04|+/-2.70E-06|Jy|2011A&A...528A..35M|uncertainty|     23.68 microns   | Broad-band measurement|12 37 09.14 +62 15 07.92 (J2000)| Flux integrated from map|                                        |From new raw data
1|MIPS 24 microns      | 128.    |+/-6.0 |microJy         |1.25E+13 |  128.E-06|+/-6.0E-06 |Jy |1990IRASF.C...0000M|3sigma uncertainty| 25        microns   | Broad-band measurement|115813.1 +302058 (B1950)| Flux in fixed aperture|                                        |From new raw data
22|70 microns (MIPS)   ||<3.0       |milliJy             |4.20E+12||3.00E-03|Jy|2011A&A...528A..35M|no uncertainty reported|     71.42 microns   | Broad-band measurement|12 37 09.14 +62 15 07.92 (J2000)| Flux integrated from map|                                        |From new raw data
2|70 microns (PACS)    |         |<2.0   |mJy             |4.283e+12|          |2.0E-03    |Jy |2.40e+01 |3sigma |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
3|100 microns (PACS)   | 2.1     |+/-0.4 |mJy             |2.998e+12|  2.1E-03 |+/-0.4E-03 |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
4|160 microns (PACS)   | 3.0     |+/-1.3 |mJy             |1.874e+12|  3.0E-03 |+/-1.3E-03 |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
5|250 microns (SPIRE)  | 8.0     |+/-2.5 |mJy             |1.199e+12|  8.0E-03 |+/-2.5e-03 |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
6|350 microns (SPIRE)  |         |<9.0   |mJy             |8.565e+11|          |9.0e-03    |Jy |2.40e+01 |3sigma |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
7|500 microns (SPIRE)  |         |<12.0  |mJy             |5.996e+11|          |12.0e-03   |Jy |2.40e+01 |3sigma |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
8|1160 microns (Penner)|         |<1.6   |mJy             |2.58442E+11|        |1.6E-03    |Jy |2004MNRAS.354..779G|3sigma uncertainty|      1200 microns   | Broad-band measurement|16 36 55.9 +40 59 12 (J2000)| Flux integrated from map|S/N = 3.66                              |From new raw data
