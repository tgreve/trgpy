
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-04-05T08:15:36PDT



Photometric Data for BzK 04171

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|3.6 microns (IRAC)  | 24.00     |+/-1.20 |microJy             |8.44E+13|  2.40E-05|+/-1.20E-06|Jy|2011AJ....141....1T|rms uncertainty|     3.550 microns   | Broad-band measurement|189.110626 62.143169 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
2|4.5 microns (IRAC)  | 27.90     |+/-1.40 |microJy             |6.67E+13|  2.79E-05|+/-1.40E-06|Jy|2011AJ....141....1T|rms uncertainty|     4.493 microns   | Broad-band measurement|189.110626 62.143169 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
3|5.8 microns (IRAC)  | 23.10     |+/-1.24 |microJy             |5.23E+13|  2.31E-05|+/-1.24E-06|Jy|2011AJ....141....1T|rms uncertainty|     5.731 microns   | Broad-band measurement|189.110626 62.143169 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
4|8.0 microns (IRAC)  | 22.00     |+/-1.23 |microJy             |3.81E+13|  2.20E-05|+/-1.23E-06|Jy|2011AJ....141....1T|rms uncertainty|     7.872 microns   | Broad-band measurement|189.110626 62.143169 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
5|16 microns (IRS)    | 125.2     |+/-15.0 |microJy             |1.90E+13|  1.25E-04|+/-1.50E-05|Jy|2011AJ....141....1T|rms uncertainty|      15.8 microns   | Broad-band measurement|189.110626 62.143169 (J2000)| From fitting to map|                                        |From new raw data
6|24 microns (MIPS)   | 139.0     |+/-6.4  |microJy             |1.27E+13|  1.39E-04|+/-6.40E-06|Jy|2011AJ....141....1T|rms uncertainty|     23.68 microns   | Broad-band measurement|189.110626 62.143169 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
7|24 microns (MIPS)   | 140.0     |+/-6.0  |microJy             |1.27E+13|  1.40E-04|+/-6.00E-06|Jy|2011AJ....141....1T|rms uncertainty|     23.68 microns   | Broad-band measurement|189.110626 62.143169 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
8|24 microns (MIPS)   | 94.       |+/-26   |uJy             |1.27E+13|94.0E-06|+/-26.0E-06|Jy|2009ApJ...694.1517D|1 sigma uncertainty|     23.68 microns   | Broad-band measurement|12 37 11.89 +62 22 11.8 (J2000)| Flux integrated from map|                                        |From new raw data
9|70 microns (MIPS)   |           |<2.6    |mJy             |4.20E+12|        |2.6E-03|Jy|2009ApJ...699.1610H|3sigma|     71.42 microns   | Broad-band measurement|221804.42 +002154.4 (J2000)| Flux in fixed aperture|                                        |From new raw data
10|70 microns (PACS)  |           |<3.2    |mJy             |4.283E+12|   |3.2E-03|Jy|2004MNRAS.354..779G|3sigma uncertainty|      1200 microns   | Broad-band measurement|16 36 55.9 +40 59 12 (J2000)| Flux integrated from map|S/N = 3.66                              |From new raw data
11|100 microns (PACS) | 2.9       |+/-0.3  |mJy             |2.998e+12| 2.9E-03 |+/-0.3.E-03 |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
12|160 microns (PACS) | 9.0       |+/-1.0  |mJy             |1.874e+12|  9.0E-03|+/-1.0E-03 |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
13|250 microns (SPIRE)| 14.5      |+/-2.5  |mJy             |1.199e+12|  14.5E-03 |+/-2.5e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
15|350 microns (SPIRE)|           |<9.0    |mJy             |8.565E+11|         |9.0E-03|Jy|2004MNRAS.354..779G|3sigma uncertainty|      1200 microns   | Broad-band measurement|16 36 55.9 +40 59 12 (J2000)| Flux integrated from map|S/N = 3.66                              |From new raw data
16|500 microns (SPIRE)|           |<12.0   |mJy                 |5.996E+11|         |12.0E-03|Jy|2004MNRAS.354..779G|3sigma uncertainty|      1200 microns   | Broad-band measurement|16 36 55.9 +40 59 12 (J2000)| Flux integrated from map|S/N = 3.66                              |From new raw data
16|850 microns (SCUBA) |           |<10.5    |mJy             |3.53E+11|        |10.5E-03|Jy|2005MNRAS.358..149P|3sigma uncertainty|     850   microns   | Broad-band measurement|12 37 11.7 +62 22 12 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
17|1160 microns (Penner)|           |<1.7    |mJy             |2.58442E+11|       |1.7E-03|Jy|2004MNRAS.354..779G|3sigma uncertainty|      1200 microns   | Broad-band measurement|16 36 55.9 +40 59 12 (J2000)| Flux integrated from map|S/N = 3.66                              |From new raw data
18|1200 microns (MAMBO)|           |<1.7    |mJy             |2.50E+11|        |1.7E-03|Jy|2004MNRAS.354..779G|3sigma uncertainty|      1200 microns   | Broad-band measurement|16 36 55.9 +40 59 12 (J2000)| Flux integrated from map|S/N = 3.66                              |From new raw data
19|43.0 GHz (VLA)      |           |<125  | microJy        |43.0E+09| |125.E-06|Jy|2006MNRAS.371..963B|2 sigma uncertainty|       1.4 GHz       | Broad-band measurement|16 36 55.767 +40 59 09.97 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
20|1.4 GHz (VLA)       | 41        |+/-7    | microJy            |1.40E+09|  4.10E-05|+/-7.00E-06|Jy|2006MNRAS.371..963B|1 sigma|       1.4 GHz       | Broad-band measurement|12 36 26.547 +62 08 35.39 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
21|1.4 GHz (VLA)       | 31.3      |+/-8.1  |microJy             |1.40E+09|  3.13E-05|+/-8.10E-06|Jy|2010ApJS..188..178M|uncertainty|       1.4 GHz       | Broad-band measurement|12 36 26.52 +62 08 35.3 (J2000)| Total flux; Beam filling or dilution corrected|Major=0.9"; Minor=0.0"; PA=178 deg      |From new raw data
22|1.4 GHz (VLA)       | 31.3      |+/-8.1  |microJy             |1.40E+09|  3.13E-05|+/-8.10E-06|Jy|2010ApJS..188..178M|uncertainty|       1.4 GHz       | Broad-band measurement|12 36 26.52 +62 08 35.3 (J2000)| Total flux; Beam filling or dilution corrected|Major=0.9"; Minor=0.0"; PA=178 deg      |From new raw data
23|1.4 GHz (VLA)       | 37.9      |+/-9.3    | microJy            |1.40E+09|  37.9E-06|+/-9.30E-06|Jy|2006MNRAS.371..963B|1 sigma|       1.4 GHz       | Broad-band measurement|12 36 26.547 +62 08 35.39 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
