

Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.

Photometric Data for SMM J02399-0136

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|350 microns (SABOCA) | 319.0 | 27. |milliJy      |8.56550e+11| 319.0E-3   |27.E-3 |Jy|2007MNRAS.376.1073Z|no uncertainty reported|     850   microns   | Broad-band measurement|02 39 51.9 -01 35 55 (J2000)| Flux integrated from map|S/N = 19.9                              |From reprocessed raw data
2|870 microns (LABOCA) | 127.0 | 10.0 |milliJy     |3.45E+11   | 127.0E-3   |10.0E-3 |Jy|2007MNRAS.376.1073Z|no uncertainty reported|     850   microns   | Broad-band measurement|02 39 51.9 -01 35 55 (J2000)| Flux integrated from map|S/N = 19.9                              |From reprocessed raw data
4|295GHz (ZSPEC) | 71.6 | 1.8 |milliJy             |2.95E+11   | 0.090886441|0.002174763 |Jy|2007MNRAS.376.1073Z|no uncertainty reported|     850   microns   | Broad-band measurement|02 39 51.9 -01 35 55 (J2000)| Flux integrated from map|S/N = 19.9                              |From reprocessed raw data
4|285GHz (ZSPEC) | 71.6 | 1.8 |milliJy             |2.85E+11   | 0.079682139|0.001914082 |Jy|2007MNRAS.376.1073Z|no uncertainty reported|     850   microns   | Broad-band measurement|02 39 51.9 -01 35 55 (J2000)| Flux integrated from map|S/N = 19.9                              |From reprocessed raw data
4|275GHz (ZSPEC) | 71.6 | 1.8 |milliJy             |2.75E+11   | 0.074544886|0.001590222 |Jy|2007MNRAS.376.1073Z|no uncertainty reported|     850   microns   | Broad-band measurement|02 39 51.9 -01 35 55 (J2000)| Flux integrated from map|S/N = 19.9                              |From reprocessed raw data
4|265GHz (ZSPEC) | 71.6 | 1.8 |milliJy             |2.65E+11   | 0.07052678 |0.001226077 |Jy|2007MNRAS.376.1073Z|no uncertainty reported|     850   microns   | Broad-band measurement|02 39 51.9 -01 35 55 (J2000)| Flux integrated from map|S/N = 19.9                              |From reprocessed raw data
4|255GHz (ZSPEC) | 59.1 | 1.2 |milliJy             |2.55E+11   | 0.060478875|0.001267365 |Jy|2007MNRAS.376.1073Z|no uncertainty reported|     850   microns   | Broad-band measurement|02 39 51.9 -01 35 55 (J2000)| Flux integrated from map|S/N = 19.9                              |From reprocessed raw data
4|245GHz (ZSPEC) | 53.7 | 1.9 |milliJy             |2.45E+11   | 0.05594415 |0.001213969 |Jy|2007MNRAS.376.1073Z|no uncertainty reported|     850   microns   | Broad-band measurement|02 39 51.9 -01 35 55 (J2000)| Flux integrated from map|S/N = 19.9                              |From reprocessed raw data
4|235GHz (ZSPEC) | 47.3 | 1.2 |milliJy             |2.35E+11   | 0.049143898|0.001507005 |Jy|2007MNRAS.376.1073Z|no uncertainty reported|     850   microns   | Broad-band measurement|02 39 51.9 -01 35 55 (J2000)| Flux integrated from map|S/N = 19.9                              |From reprocessed raw data
3|1300 microns (SMA) | 47.0 | 14.1 |milliJy        |2.30610E+11| 47.0E-3    |14.1E-3     |Jy|2007MNRAS.376.1073Z|no uncertainty reported|     850   microns   | Broad-band measurement|02 39 51.9 -01 35 55 (J2000)| Flux integrated from map|S/N = 19.9                              |From reprocessed raw data
4|225GHz (ZSPEC) | 45.2 | 1.2 |milliJy             |2.25E+11   | 0.04411366 |0.001252055 |Jy|2007MNRAS.376.1073Z|no uncertainty reported|     850   microns   | Broad-band measurement|02 39 51.9 -01 35 55 (J2000)| Flux integrated from map|S/N = 19.9                              |From reprocessed raw data
4|1360 microns (SPT) | 40.8 | 5.2 |milliJy         |2.20436E+11| 40.8E-3    |5.2E-3      |Jy|2007MNRAS.376.1073Z|no uncertainty reported|     850   microns   | Broad-band measurement|02 39 51.9 -01 35 55 (J2000)| Flux integrated from map|S/N = 19.9                              |From reprocessed raw data
4|215GHz (ZSPEC) | 37.2 | 1.2 |milliJy             |2.15E+11   | 0.037629954|0.001284752 |Jy|2007MNRAS.376.1073Z|no uncertainty reported|     850   microns   | Broad-band measurement|02 39 51.9 -01 35 55 (J2000)| Flux integrated from map|S/N = 19.9                              |From reprocessed raw data
4|205GHz (ZSPEC) | 34.0 | 1.8 |milliJy             |2.05E+11   | 0.034354109|0.001787242 |Jy|2007MNRAS.376.1073Z|no uncertainty reported|     850   microns   | Broad-band measurement|02 39 51.9 -01 35 55 (J2000)| Flux integrated from map|S/N = 19.9                              |From reprocessed raw data
5|2100 microns (SPT) | 13.4 | 2.0 |milliJy         |1.42758E+11| 13.4E-3    |2.0E-3      |Jy|2007MNRAS.376.1073Z|no uncertainty reported|     850   microns   | Broad-band measurement|02 39 51.9 -01 35 55 (J2000)| Flux integrated from map|S/N = 19.9                              |From reprocessed raw data
