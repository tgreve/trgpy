
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-07-10T13:42:15PDT



Photometric Data for SPT0551-50

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
3|100 microns (PACS) | 13.3      |+/-2.5  |mJy             |2.998e+12|13.3E-03|+/-2.5E-03             |Jy|2005MNRAS.358..149P|uncertainty|     850   microns   | Broad-band measurement|12 37 11.7 +62 22 12 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
4|160 microns (PACS) | 63.4     |+/-13.7 |mJy                |1.874e+12|63.4E-03|+/-13.7E-03  |Jy |2.40e+01          |3sigma|-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
5|250 microns (SPIRE)| 148.8    |+/-7.1 |mJy                 |1.199e+12| 148.8E-03|+/-7.1e-03 |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
6|350 microns (SPIRE)| 189.9    |+/-7.3  |mJy                |8.565e+11|189.9E-03 |+/-7.3e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
8|500 microns (SPIRE) | 196.9   |+/-7.5 |mJy                 |5.996e+11|196.9E-03 |+/-7.5e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
1|870 microns (LABOCA)| 74.0    |+/-6.3  |milliJy            |3.45E+11|  74.0E-03|+/-6.3E-03|Jy|2009ApJ...707.1201W|uncertainty|       870 microns   | Broad-band measurement|03 32 29.33 -27 56 19.3 (J2000)| Flux integrated from map|S/N = 4.6                               |From new raw data
1|1.4 mm (SPT)        | 27.0    |+/-4.2 |milliJy             |2.20E+11|  27.0E-03|+/-4.2E-03|Jy|2010ApJ...719..763V|uncertainty|       1.4 mm        | Broad-band measurement|74.804 -59.708 (J2000)| Flux integrated from map|De-boosted flux; S/N = 7.05             |From new raw data
3|2.0 mm (SPT)        | 5.0     |+/-0.9 |milliJy             |1.50E+11|  5.0E-03|+/-0.9E-03|Jy|2010ApJ...719..763V|uncertainty|       2.0 mm        | Broad-band measurement|74.804 -59.708 (J2000)| Flux integrated from map|De-boosted flux; S/N = 6.20             |From new raw data
3|3.0 mm (SPT)        | 1.04    |+/-0.17 |milliJy            |9.99E+10|  1.04E-03|+/-0.17E-03|Jy|2010ApJ...719..763V|uncertainty|       2.0 mm        | Broad-band measurement|74.804 -59.708 (J2000)| Flux integrated from map|De-boosted flux; S/N = 6.20             |From new raw data
