
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-02-19T11:57:36PST



Photometric Data for SMM J13120+4242

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|H{beta} (Keck)      | 0.18E-16  |+/-0.15E-16|ergs cm^-2^ s^-1^   |6.17E+14|  2.92E-09|+/-2.43E-09|Jy|2006ApJ...651..713T|uncertainty|    4861   A         | Line measurement; flux integrated over line; lines measured in emission| | Flux integrated from map|                                        |From new raw data
2|[O III] 4959 (Keck) | 0.27E-16  |+/-0.19E-16|ergs cm^-2^ s^-1^   |6.05E+14|  4.46E-09|+/-3.14E-09|Jy|2006ApJ...651..713T|uncertainty|    4959   A         | Line measurement; flux integrated over line; lines measured in emission| | Flux integrated from map|                                        |From new raw data
3|[O III] 5007 (Keck) | 0.79E-16  |+/-0.19E-16|ergs cm^-2^ s^-1^   |5.99E+14|  1.32E-08|+/-3.17E-09|Jy|2006ApJ...651..713T|uncertainty|    5007   A         | Line measurement; flux integrated over line; lines measured in emission| | Flux integrated from map|                                        |From new raw data
4|R (SUBARU)          | 24.2      |+/-0.3  |mag                 |4.76E+14|  6.52E-07|+/-1.80E-07|Jy|2006ApJS..167..103F|rms uncertainty|    6300   A         | Broad-band measurement| | Flux in fixed aperture|3" radius aperture                      |From new raw data
5|I (Cousins)         | 23.10     |+/-0.06 |mag                 |3.79E+14|  1.47E-06|+/-8.34E-08|Jy|2004ApJ...616...71S|1 sigma|    7900   A         | Broad-band measurement| | Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
6|z (SUBARU)          | 23.0      |+/-0.5  |mag                 |3.26E+14|  1.38E-06|+/-6.36E-07|Jy|2006ApJS..167..103F|rms uncertainty|    9200   A         | Broad-band measurement| | Flux in fixed aperture|3" radius aperture                      |From new raw data
7|J (2MASS)           | 22.18     |+/-0.26 |mag                 |2.40E+14|  2.14E-06|+/-5.78E-07|Jy|2004ApJ...616...71S|1 sigma|    1.25   microns   | Broad-band measurement| | Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
8|F160W (HST) AB      | 22.87     |+/-0.08 |mag                 |1.87E+14|  2.58E-06|+/-1.90E-07|Jy|2010MNRAS.405..234S|uncertainty|      1.60 microns   | Broad-band measurement|13 12 01.17 +42 42 08.1 (J2000)| Flux in fixed aperture|                                        |From new raw data
9|K_s_ (2MASS)        | 20.47     |+/-0.21 |mag                 |1.38E+14|  4.33E-06|+/-9.23E-07|Jy|2004ApJ...616...71S|1 sigma|    2.17   microns   | Broad-band measurement| | Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
10|3.6 microns (IRAC)  | 10.9      |+/-1.3  |microJy             |8.44E+13|  1.09E-05|+/-1.30E-06|Jy|2009ApJ...699.1610H|uncertainty|     3.550 microns   | Broad-band measurement|13 12 01.18 +42 42 08.3 (J2000)| Flux in fixed aperture|                                        |From new raw data
11|4.5 microns (IRAC)  | 15.5      |+/-2.0  |microJy             |6.67E+13|  1.55E-05|+/-2.00E-06|Jy|2009ApJ...699.1610H|uncertainty|     4.493 microns   | Broad-band measurement|13 12 01.18 +42 42 08.3 (J2000)| Flux in fixed aperture|                                        |From new raw data
12|5.8 microns (IRAC)  | 24.8      |+/-3.8  |microJy             |5.23E+13|  2.48E-05|+/-3.80E-06|Jy|2009ApJ...699.1610H|uncertainty|     5.731 microns   | Broad-band measurement|13 12 01.18 +42 42 08.3 (J2000)| Flux in fixed aperture|                                        |From new raw data
13|8.0 microns (IRAC)  | 30.2      |+/-4.2  |microJy             |3.85E+13|  3.02E-05|+/-4.20E-06|Jy|2009ApJ...699.1610H|uncertainty|     7.782 microns   | Broad-band measurement|13 12 01.18 +42 42 08.3 (J2000)| Flux in fixed aperture|                                        |From new raw data
14|350 microns (SHARC2)| 21.1      |+/-7.7  |milliJy             |8.57E+11|  2.11E-02|+/-7.70E-03|Jy|2006ApJ...650..592K|uncertainty|     350   microns   | Broad-band measurement| | Total flux|                                        |From new raw data
15|CO(6-5) (PdBI)      | 2.54      |+/-0.1  |Jy km/s             |6.91E+11|  4.36E-07|+/-1.72E-08|Jy|2010ApJ...724..233E|uncertainty|   691.473 GHz       | Line measurement; flux integrated over line; lines measured in emission| | Flux integrated from map|                                        |From new raw data
16|CO(4-3) line (IRAM) | 1.7       |+/-0.3  |Jy km s^-1^         |4.61E+11|  2.92E-07|+/-5.15E-08|Jy|2005MNRAS.359.1165G|uncertainty|   3.408             | Line measurement; flux integrated over line; lines measured in emission|13 12 01.20 +42 42 08.8 (J2000)| Flux integrated from map|                                        |From new raw data
17|850 microns (SCUBA) | 6.2       |+/-1.2  |milliJy             |3.53E+11|  6.20E-03|+/-1.20E-03|Jy|2005ApJ...622..772C|uncertainty|     850   microns   | Broad-band measurement|131201.17 +424208.1 (J2000)| Flux integrated from map|                                        |From new raw data
18|2.6mm  (pdbi)       |           |<60     |microJy             |1.15E+11|  |60.E-06|Jy|2006ApJ...650..592K|3sigma uncertainty|     350   microns   | Broad-band measurement| | Total flux|                                        |From new raw data
19|1.4 GHz (VLA)       | 59        |+/-16   |microJy             |1.40E+09|  5.90E-05|+/-1.60E-05|Jy|2006ApJS..167..103F|uncertainty|     1.4   GHz       | Broad-band measurement|13 12 01.172 +42 42 08.39 (J2000)| Flux integrated from map|Corrected to the sky; see paper         |From new raw data
