

Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.


queryDateTime:2009-11-03T15:07:35PST






Photometric Data for MIPS16144 (z=2.131)

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
0|R (Cousins)         | 23.3     |+/-0.2  |mag                 |4.72E+14|  1.73781e-06|+/-3.51490e-07 |Jy|2004ApJ...616...71S|sigma uncertainty|    1.25   microns   | Broad-band measurement| | Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
1|R (KPNO)            | 1.692     ||microJy             |4.66E+14|  1.69E-06||Jy|2007ApJ...658..778Y|no uncertainty reported|    6440   A         | Broad-band measurement|172422.10 +593150.8 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data
2|R (Cousins) m_tot   | 23.10     |+/-0.08 |mag                 |4.65E+14|  1.76E-06|+/-1.30E-07|Jy|2004AJ....128....1F|based on count statistics only|6440       A         | Broad-band measurement|172421.911 +593151.27 (J2000)| Total flux|                                        |From new raw data
3|R (Cousins) m_aper  | 23.45     |+/-0.07 |mag                 |4.65E+14|  1.28E-06|+/-8.22E-08|Jy|2004AJ....128....1F|based on count statistics only|6440       A         | Broad-band measurement|172421.911 +593151.27 (J2000)| Flux in fixed aperture|3-arcsecond aperture                    |From new raw data
4|F160W (HST NICMOS)         | 20.36     ||mag                 |1.87E+14|  7.49E-06||Jy|2011ApJ...730..125Z|no uncertainty reported|      1.60 microns   | Broad-band measurement|| Flux integrated from map|                                        |From new raw data
5|F160W (HST NICMOS)         | 20.85     || mag                |1.86E+14|  4.77E-06||Jy|2008ApJ...680..232D|no uncertainty reported|      1.61 microns   | Broad-band measurement|17 24 22.03 +59 31 50.63 (J2000)| Flux integrated from map|                                        |From new raw data
6|3.6 microns (IRAC)  | 68        |+/-3    | microJy            |8.44E+13|  6.80E-05|+/-3.00E-06|Jy|2007ApJ...664..713S|uncertainty|   3.550   microns   | Broad-band measurement|| Flux in fixed aperture|7.3" diameter aperture                  |From reprocessed raw data
7|3.6 microns (IRAC)  | 65.75     |+/-7.55 |microJy             |8.42E+13|  6.57E-05|+/-7.55E-06|Jy|2005ApJS..161...41L|uncertainty|3.56       microns   | Broad-band measurement|172422.03 +593150.6 (J2000)| Flux in fixed aperture|Aperture =       7.59 arcsec.           |From new raw data
8|4.5 microns (IRAC)  | 84        |+/-3    | microJy            |6.67E+13|  8.40E-05|+/-3.00E-06|Jy|2007ApJ...664..713S|uncertainty|   4.493   microns   | Broad-band measurement|| Flux in fixed aperture|7.3" diameter aperture                  |From reprocessed raw data
9|4.5 microns (IRAC)  | 87.84     |+/-9.76 |microJy             |6.63E+13|  8.78E-05|+/-9.76E-06|Jy|2005ApJS..161...41L|uncertainty|4.52       microns   | Broad-band measurement|172422.03 +593150.6 (J2000)| Flux in fixed aperture|Aperture =       7.59 arcsec.           |From new raw data
10|5.8 microns (IRAC)  | 108       |+/-24   | microJy            |5.23E+13|  1.08E-04|+/-2.40E-05|Jy|2007ApJ...664..713S|uncertainty|   5.731   microns   | Broad-band measurement|| Flux in fixed aperture|7.3" diameter aperture                  |From reprocessed raw data
11|5.8 microns (IRAC)  | 119.79    |+/-20.16|microJy             |5.23E+13|  1.20E-04|+/-2.02E-05|Jy|2005ApJS..161...41L|uncertainty|5.73       microns   | Broad-band measurement|172422.03 +593150.6 (J2000)| Flux in fixed aperture|Aperture =       7.59 arcsec.           |From new raw data
14|8.0 microns (IRAC)  | 94.712    ||microJy             |3.81E+13|  9.47E-05||Jy|2007ApJ...658..778Y|no uncertainty reported|   7.872   microns   | Broad-band measurement|172422.10 +593150.8 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data
15|8.0 microns (IRAC)  | 105       |+/-19   | microJy            |3.81E+13|  1.05E-04|+/-1.90E-05|Jy|2007ApJ...664..713S|uncertainty|   7.872   microns   | Broad-band measurement|| Flux in fixed aperture|7.3" diameter aperture                  |From reprocessed raw data
16|8.0 microns (IRAC)  | 108.24    |+/-15.96|microJy             |3.79E+13|  1.08E-04|+/-1.60E-05|Jy|2005ApJS..161...41L|uncertainty|7.91       microns   | Broad-band measurement|172422.03 +593150.6 (J2000)| Flux in fixed aperture|Aperture =       7.59 arcsec.           |From new raw data
17|8 microns (IRAC) | 1.8       |+/-1   %|milliJy             |3.75E+13|  1.80E-03|+/-1.80E-05|Jy|2009ApJ...698.1682W|typical accuracy|         8 microns   | Broad-band measurement|17 24 22.10 +59 31 50.8 (J2000)| Peak flux|                                        |From reprocessed raw data
20|24 microns (MIPS)   | 1010.148  ||microJy             |1.27E+13|  1.01E-03||Jy|2007ApJ...658..778Y|no uncertainty reported|   23.68   microns   | Broad-band measurement|172422.10 +593150.8 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data; measurementmodified from published value
1|MIPS 24um           | 1.12     |+/-0.3  |milliJy             |1.27E+13|  1.12E-03|+/-0.34E-03 |Jy|1996AJ....111.1431B|uncertainty|1.49       GHz       | Broad-band measurement| | Peak flux|                                        |From new raw data
2|MIPS 70um           |          |<3.6    |milliJy             |4.20E+12|          |4.6E-03|Jy|2010Natur.464..733S|3sigma uncertainty|     71.42 microns   | Broad-band measurement|21 35 11.6 -01 02 52.0 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
21|70 microns (MIPS)   | 2.2       |+/-1.2  | milliJy            |4.20E+12|  2.20E-03|+/-1.20E-03|Jy|2007ApJ...664..713S|estimated error|   71.42   microns   | Broad-band measurement|| Flux in fixed aperture|3 pixel radius aperture                 |From reprocessed raw data
3|MIPS 160um          |          |<30     |milliJy             |1.92E+12|          |30.0E-03|Jy|2009A&A...502..541E|3 sigma|     155.9 microns   | Broad-band measurement| | Flux in fixed aperture|                                        |From reprocessed raw data
4|MAMBO 1200um        | 2.93     |+/-0.59 |milliJy             |2.50E+11|  2.93E-03|+/-0.59E-03|Jy|2004MNRAS.354..779G|uncertainty|      1200 microns   | Broad-band measurement|16 37 06.7 +40 53 15 (J2000)| Flux integrated from map|S/N = 3.81                              |From new raw data
5|PDBI 2.7mm MONO     | 0.5      |+/-0.1 |milliJy             |1.10E+11|  0.5E-03|+/-0.1E-03|Jy|2004MNRAS.354..779G|uncertainty|      1200 microns   | Broad-band measurement|16 37 06.7 +40 53 15 (J2000)| Flux integrated from map|S/N = 3.81                              |From new raw data
6|VLA 1.4GHz          | 0.12     |+/-0.03 |milliJy             |1.4E9   |  0.12E-3 |+/-0.03E-3|Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
