
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-06-17T13:31:37PDT



Photometric Data for GOODS J123702.71+621426.6

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|U_n AB              | 28.13     |+/-0.72 |mag                 |8.44E+14|  2.03E-08|+/-1.35E-08|Jy|2003ApJ...592..728S|typical accuracy|    3550   A         | Broad-band measurement|12 37 02.70 +62 14 26.3 (J2000)| Flux in fixed aperture|2" diameter aperture                    |From new raw data; derived from a flux in a different bandand a color
2|U (KPNO) AB         | 28.13     ||mag                 |8.44E+14|  2.03E-08||Jy|2006ApJ...653.1004R|no uncertainty reported|    3550   A         | Broad-band measurement|123702.68 +621425.9 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data; derived from aflux in a different band and a color
3|U (KPNO) AB         | 26.4      || mag                |8.22E+14|  1.00E-07||Jy|2004AJ....127.3137C|no uncertainty reported| 3647.65   A         | Broad-band measurement|189.261368 +62.24059 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
4|B (Subaru) AB       | 25.2      || mag                |6.77E+14|  3.02E-07||Jy|2004AJ....127.3137C|no uncertainty reported| 4427.60   A         | Broad-band measurement|189.261368 +62.24059 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
5|G (KECK) AB         | 25.70     ||mag                 |6.27E+14|  1.91E-07||Jy|2006ApJ...653.1004R|no uncertainty reported|    4780   A         | Broad-band measurement|123702.68 +621425.9 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data; derived from aflux in a different band and a color
6|G AB                | 25.70     |+/-0.18 |mag                 |6.27E+14|  1.91E-07|+/-3.16E-08|Jy|2003ApJ...592..728S|typical accuracy|    4780   A         | Broad-band measurement|12 37 02.70 +62 14 26.3 (J2000)| Flux in fixed aperture|2" diameter aperture                    |From new raw data; derived from a flux in a different bandand a color
7|V (Subaru) AB       | 24.6      || mag                |5.48E+14|  5.25E-07||Jy|2004AJ....127.3137C|no uncertainty reported| 5471.22   A         | Broad-band measurement|189.261368 +62.24059 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
8|R (Keck II) AB      | 24.46     || mag                |4.62E+14|  5.97E-07||Jy|2004AJ....127.3121W|no uncertainty reported|   648.7   A         | Broad-band measurement|12 37 02.709 +62 14 26.21 (J2000)| Total flux|                                        |From new raw data
9|R (Subaru) AB       | 24.2      || mag                |4.59E+14|  7.59E-07||Jy|2004AJ....127.3137C|no uncertainty reported| 6534.16   A         | Broad-band measurement|189.261368 +62.24059 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
10|R (KECK) AB         | 24.61     ||mag                 |4.39E+14|  5.20E-07||Jy|2006ApJ...653.1004R|no uncertainty reported|    6830   A         | Broad-band measurement|123702.68 +621425.9 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data
11|R AB                | 24.61     |+/-0.1  |mag                 |4.39E+14|  5.20E-07|+/-4.79E-08|Jy|2003ApJ...592..728S|typical accuracy|    6830   A         | Broad-band measurement|12 37 02.70 +62 14 26.3 (J2000)| Total flux|                                        |From new raw data
12|I (Subaru) AB       | 24.0      || mag                |3.76E+14|  9.12E-07||Jy|2004AJ....127.3137C|no uncertainty reported| 7975.89   A         | Broad-band measurement|189.261368 +62.24059 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
13|z' (Subaru) AB      | 23.9      || mag                |3.31E+14|  1.00E-06||Jy|2004AJ....127.3137C|no uncertainty reported| 9069.21   A         | Broad-band measurement|189.261368 +62.24059 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
14|HK' (UH) AB         | 22.0      || mag                |1.58E+14|  5.75E-06||Jy|2004AJ....127.3137C|no uncertainty reported|18947.38   A         | Broad-band measurement|189.261368 +62.24059 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
15|3.6 microns IRAC AB | 20.83     |+/-0.07 |mag                 |8.44E+13|  1.69E-05|+/-1.09E-06|Jy|2006ApJ...653.1004R|uncertainty|   3.550   microns   | Broad-band measurement|123702.68 +621425.9 (J2000)| Flux integrated from map|                                        |From new raw data
16|3.6 microns IRAC AB | 21.01     |+/-0.09 |mag                 |8.44E+13|  1.43E-05|+/-1.19E-06|Jy|2010MNRAS.401.1521M|uncertainty|     3.550 microns   | Broad-band measurement|| Total flux|                                        |Averaged from previously published data
17|4.5 microns IRAC AB | 20.88     |+/-0.07 |mag                 |6.67E+13|  1.61E-05|+/-1.04E-06|Jy|2006ApJ...653.1004R|uncertainty|   4.493   microns   | Broad-band measurement|123702.68 +621425.9 (J2000)| Flux integrated from map|                                        |From new raw data
18|4.5 microns IRAC AB | 21.16     |+/-0.07 |mag                 |6.67E+13|  1.25E-05|+/-8.04E-07|Jy|2010MNRAS.401.1521M|uncertainty|     4.493 microns   | Broad-band measurement|| Total flux|                                        |Averaged from previously published data
19|5.8 microns IRAC AB | 21.04     |+/-0.07 |mag                 |5.23E+13|  1.39E-05|+/-8.98E-07|Jy|2006ApJ...653.1004R|uncertainty|   5.731   microns   | Broad-band measurement|123702.68 +621425.9 (J2000)| Flux integrated from map|                                        |From new raw data
20|5.8 microns IRAC AB | 21.08     |+/-0.07 |mag                 |5.23E+13|  1.34E-05|+/-8.66E-07|Jy|2010MNRAS.401.1521M|uncertainty|     5.731 microns   | Broad-band measurement|| Total flux|                                        |Averaged from previously published data
21|8.0 microns IRAC AB | 21.08     |+/-0.07 |mag                 |3.81E+13|  1.34E-05|+/-8.66E-07|Jy|2006ApJ...653.1004R|uncertainty|   7.872   microns   | Broad-band measurement|123702.68 +621425.9 (J2000)| Flux integrated from map|                                        |From new raw data
22|8.0 microns IRAC AB | 21.10     |+/-0.07 |mag                 |3.81E+13|  1.32E-05|+/-8.50E-07|Jy|2010MNRAS.401.1521M|uncertainty|     7.872 microns   | Broad-band measurement|| Total flux|                                        |Averaged from previously published data
23|24 microns (MIPS)   | 26.4      |+/-3.0  |microJy             |1.27E+13|  2.64E-05|+/-3.00E-06|Jy|2011A&A...528A..35M|uncertainty|     23.68 microns   | Broad-band measurement|12 37 02.70 +62 14 26.08 (J2000)| Flux integrated from map|                                        |From new raw data
24|70 microns (MIPS)   ||<2.7       |milliJy             |4.20E+12||2.70E-03|Jy|2011A&A...528A..35M|no uncertainty reported|     71.42 microns   | Broad-band measurement|12 37 02.70 +62 14 26.08 (J2000)| Flux integrated from map|                                        |From new raw data
25|1.4 GHz (VLA)       | 21.5      |+/-4.2  |microJy             |1.40E+09|  2.15E-05|+/-4.20E-06|Jy|2010ApJS..188..178M|uncertainty|       1.4 GHz       | Broad-band measurement|12 37 02.57 +62 14 26.6 (J2000)| Total flux; Beam filling or dilution corrected|Major=0.0"; Minor=0.0"; PA=0 deg        |From new raw data
