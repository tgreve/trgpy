

Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.


queryDateTime:2009-11-03T15:07:35PST






Photometric Data for MIPS429 (z=2.201)

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|R (Cousins) AB      |           |<25.71  |mag                   |4.72E+14|          |1.888e-07|Jy|2004ApJ...616...71S|3sigma uncertainty|    1.25   microns   | Broad-band measurement| | Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
1|R (KPNO)            | 0.560     ||microJy             |4.66E+14|  5.60E-07||Jy|2007ApJ...658..778Y|no uncertainty reported|    6440   A         | Broad-band measurement|171611.81 +591213.3 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data
2|R (Cousins) m_tot   | 24.30     |+/-0.20 |mag                 |4.65E+14|  5.83E-07|+/-1.07E-07|Jy|2004AJ....128....1F|based on count statistics only|6440       A         | Broad-band measurement|171611.807 +591213.53 (J2000)| Total flux|                                        |From new raw data
3|R (Cousins) m_aper  | 24.58     |+/-0.16 |mag                 |4.65E+14|  4.51E-07|+/-6.64E-08|Jy|2004AJ....128....1F|based on count statistics only|6440       A         | Broad-band measurement|171611.807 +591213.53 (J2000)| Flux in fixed aperture|3-arcsecond aperture                    |From new raw data
4|3.6 microns (IRAC)  | 18        |+/-6    | microJy            |8.44E+13|  1.80E-05|+/-6.00E-06|Jy|2007ApJ...664..713S|uncertainty|   3.550   microns   | Broad-band measurement|| Flux in fixed aperture|7.3" diameter aperture                  |From reprocessed raw data
5|4.5 microns (IRAC)  | 6         |+/-4    | microJy            |6.67E+13|  6.00E-06|+/-4.00E-06|Jy|2007ApJ...664..713S|uncertainty|   4.493   microns   | Broad-band measurement|| Flux in fixed aperture|7.3" diameter aperture                  |From reprocessed raw data
6|5.8 microns (IRAC)  | 4         |+/-24   | microJy            |5.23E+13|  4.00E-06|+/-2.40E-05|Jy|2007ApJ...664..713S|uncertainty|   5.731   microns   | Broad-band measurement|| Flux in fixed aperture|7.3" diameter aperture                  |From reprocessed raw data
10|8.0 microns (IRAC)  | 20.000    ||microJy             |3.81E+13|  2.00E-05||Jy|2007ApJ...658..778Y|no uncertainty reported|   7.872   microns   | Broad-band measurement|171611.81 +591213.3 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data
11|8 microns (IRAC) | 1.4       |+/-1   %|milliJy             |3.75E+13|  1.40E-03|+/-1.40E-05|Jy|2009ApJ...698.1682W|typical accuracy|         8 microns   | Broad-band measurement|17 16 11.81 +59 12 13.3 (J2000)| Peak flux|                                        |From reprocessed raw data
1|MIPS 24um           | 1.10     |+/-0.33 |milliJy             |1.27E+13|  1.10E-03|+/-0.33E-03 |Jy|1996AJ....111.1431B|uncertainty|1.49       GHz       | Broad-band measurement| | Peak flux|                                        |From new raw data
13|24 microns (MIPS)   | 1.10      |+/-0.06 |milliJy             |1.27E+13|  1.10E-03|+/-6.00E-05|Jy|2006AJ....131.2859F|uncertainty|   23.68   microns   | Broad-band measurement|171611.842 +591213.16 (J2000)| From fitting to map|S/N = 17.1                              |From new raw data
2|MIPS 70um           |          |<4.5    |milliJy             |4.20E+12|          |4.5E-03|Jy|2010Natur.464..733S|3 sigma|     71.42 microns   | Broad-band measurement|21 35 11.6 -01 02 52.0 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
15|70 microns (MIPS)   | 3.5       |+/-1.5  | milliJy            |4.20E+12|  3.50E-03|+/-1.50E-03|Jy|2007ApJ...664..713S|estimated error|   71.42   microns   | Broad-band measurement|| Flux in fixed aperture|3 pixel radius aperture                 |From reprocessed raw data
3|MIPS 160um          |          |<30     |milliJy             |1.92E+12|          |30.0E-03|Jy|2009A&A...502..541E|3 sigma|     155.9 microns   | Broad-band measurement| | Flux in fixed aperture|                                        |From reprocessed raw data
4|MAMBO 1200um        | 1.03     |+/-0.57 |milliJy             |2.50E+11|  1.03E-03|+/-0.57E-03|Jy|2004MNRAS.354..779G|uncertainty|      1200 microns   | Broad-band measurement|16 37 06.7 +40 53 15 (J2000)| Flux integrated from map|S/N = 3.81                              |From new raw data
5|VLA 1.4GHz          |          |<0.08   |milliJy             |1.4E+09 |          |0.08E-3 |Jy |2003MNRAS.343..293M|3sigma uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
