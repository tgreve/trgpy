
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-06-17T16:55:06PDT



Photometric Data for 4C +60.07

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|0.5-8 keV (Chandra) | 8.2E-15   |+/-1.6E-15|erg/s/cm^2^         |1.03E+18|  7.96E-10|+/-1.55E-10|Jy|2009ApJ...702L.114S|uncertainty|     4.25  keV       | Broad-band measurement|| Modelled datum|                                        |From new raw data; Extinction-corrected for Milky Way; NEDfrequency assigned to mid-point of band in keV
2|3.6 microns (IRAC)  | 27.3      |+/-3.1  | microJy            |8.44E+13|  2.73E-05|+/-3.10E-06|Jy|2007ApJS..171..353S|uncertainty|   3.550   microns   | Broad-band measurement|05 12 54.8 +60 30 52.01 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
3|4.5 microns (IRAC)  | 33.6      |+/-3.7  | microJy            |6.67E+13|  3.36E-05|+/-3.70E-06|Jy|2007ApJS..171..353S|uncertainty|   4.493   microns   | Broad-band measurement|05 12 54.8 +60 30 52.01 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
4|5.8 microns (IRAC)  | 35.1      |+/-8.4  | microJy            |5.23E+13|  3.51E-05|+/-8.40E-06|Jy|2007ApJS..171..353S|uncertainty|   5.731   microns   | Broad-band measurement|05 12 54.8 +60 30 52.01 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
5|8.0 microns (IRAC)  | 37.2      |+/-9.5  | microJy            |3.81E+13|  3.72E-05|+/-9.50E-06|Jy|2007ApJS..171..353S|uncertainty|   7.872   microns   | Broad-band measurement|05 12 54.8 +60 30 52.01 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
6|16 microns (IRS)    | 175.0     |+/-33.0 | microJy            |1.87E+13|  1.75E-04|+/-3.30E-05|Jy|2007ApJS..171..353S|uncertainty|      16   microns   | Broad-band measurement|05 12 54.8 +60 30 52.01 (J2000)| Flux in fixed aperture|6" diameter aperture                    |From reprocessed raw data
7|24 microns (MIPS)   | 1340.0    |+/-83.7 | microJy            |1.27E+13|  1.34E-03|+/-8.37E-05|Jy|2007ApJS..171..353S|uncertainty|   23.68   microns   | Broad-band measurement|05 12 54.8 +60 30 52.01 (J2000)| Flux in fixed aperture|13" diameter aperture                   |From reprocessed raw data
8|70 microns (MIPS)   ||<3750      | microJy            |4.20E+12||3.75E-03|Jy|2007ApJS..171..353S|3 sigma|   71.42   microns   | Broad-band measurement|05 12 54.8 +60 30 52.01 (J2000)| Flux in fixed aperture|35" diameter aperture                   |From reprocessed raw data
9|160 microns (MIPS)  ||<64600     | microJy            |1.92E+12||6.46E-02|Jy|2007ApJS..171..353S|3 sigma|   155.9   microns   | Broad-band measurement|05 12 54.8 +60 30 52.01 (J2000)| Flux in fixed aperture|50" diameter aperture                   |From reprocessed raw data
10|450 microns (SCUBA) | 10        |+/-13   | milliJy            |6.66E+11|  1.00E-02|+/-1.30E-02|Jy|2004MNRAS.353..377R|uncertainty|       450 microns   | Broad-band measurement|05 12 55.15 +60 30 51.0 (J2000)| Not reported in paper|Good quality data                       |From new raw data
11|850 microns (SCUBA) | 17        |+/-1    |milliJy             |3.53E+11|  1.70E-02|+/-1.00E-03|Jy|2007MNRAS.375.1299V|uncertainty|     850   microns   | Broad-band measurement|| Flux integrated from map|From 2001MNRAS.323..417A                |Averaged from previously published data
12|850 microns (SCUBA) | 11.5      |+/-1.5  | milliJy            |3.53E+11|  1.15E-02|+/-1.50E-03|Jy|2004MNRAS.353..377R|uncertainty|       850 microns   | Broad-band measurement|05 12 55.15 +60 30 51.0 (J2000)| Not reported in paper|Good quality data                       |From new raw data
13|CO (1-0) (VLA)      | 0.09      |+/-0.01 | Jy km/s            |1.15E+11|  7.23E+03|+/-8.03E+02|Jy-Hz|2004A&A...419...99G|uncertainty|   3.788             | Line measurement; flux integrated over line; lines measured in emission|05 12 55.30 +60 30 52.29 (J2000)| Flux integrated from map|Narrow component                        |From new raw data
14|CO (1-0) (VLA)      | 0.15      |+/-0.03 | Jy km/s            |1.15E+11|  1.20E+04|+/-2.41E+03|Jy-Hz|2004A&A...419...99G|uncertainty|   3.788             | Line measurement; flux integrated over line; lines measured in emission|05 12 54.75 +60 30 50.92 (J2000)| Flux integrated from map|Broad component                         |From new raw data
15|1.4GHz              | 156.8     |+/-4.7  |milliJy             |1.40E+09|  1.57E-01|+/-4.70E-03|Jy|1998AJ....115.1693C|uncertainty|    1.40   GHz       | Broad-band measurement|05 12 54.86 +60 30 52.0 (J2000)| Flux integrated from map|                                        |From new raw data
16|365 MHz (Texas)     | 1.242     |+/-0.041|Jy                  |3.65E+08|  1.24E+00|+/-4.10E-02|Jy|1996AJ....111.1945D|internal error|365        MHz       | Broad-band measurement; obtained by interpolation over frequency|050826.064 602718.85 (B1950)| Integrated from scans|Model:P;MFlag:+;EFlag:+;LFlag:+.        |From new raw data
17|178 MHz             | 3.1       |+/-15.0%|Jy                  |1.78E+08|  3.10E+00|+/-4.65E-01|Jy|1967MmRAS..71...49G|uncertainty|178        MHz       | Broad-band measurement|050825.5 +602642 (B1950)| Integrated from scans|                                        |From new raw data; Uncorrected for known sources in beam
18|151 MHz (6C)        | 3.47      |+/-0.130|Jy                  |1.52E+08|  3.47E+00|+/-1.30E-01|Jy|1993MNRAS.262.1057H|typical accuracy|151.5      MHz       | Broad-band measurement|050826.0 602714. (B1950)| Flux integrated from map|                                        |From new raw data
19|151 MHz (6C)        | 3.50      |+/-0.060|Jy                  |1.52E+08|  3.50E+00|+/-6.00E-02|Jy|1993MNRAS.262.1057H|typical accuracy|151.5      MHz       | Broad-band measurement|050826.0 602714. (B1950)| Peak flux|                                        |From new raw data
20|74 MHz (VLA)        | 8.93      |+/-0.92 | Jy                 |7.38E+07|  8.93E+00|+/-9.20E-01|Jy|2007AJ....134.1245C|rms uncertainty|    73.8   MHz       | Broad-band measurement|05 12 54.98 +60 30 53.1 (J2000)| Flux integrated from map|Corrected for clean bias                |From new raw data
21|38 MHz (8C)         | 15.6      |+/-10.0%|Jy                  |3.78E+07|  1.56E+01|+/-1.56E+00|Jy|1995MNRAS.274..447H|no uncertainty reported|38         MHz       | Broad-band measurement|050827. +602656. (B1950)| Flux integrated from map|Single component source                 |From new raw data
22|38 MHz (8C)         | 12.7      |+/-10.0%|Jy                  |3.78E+07|  1.27E+01|+/-1.27E+00|Jy|1995MNRAS.274..447H|no uncertainty reported|38         MHz       | Broad-band measurement|050827. +602656. (B1950)| Peak flux|Single component source                 |From new raw data
