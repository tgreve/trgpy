
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-07-10T07:30:04PDT



Photometric Data for 2MASSi J1612399+471157

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|u (SDSS PSF) AB     | 17.738    |+/-0.026|asinh mag           |8.36E+14|  3.03E-04|+/-7.25E-06|Jy|2007SDSS6.C...0000:|based on count statistics only|3585       A         | Broad-band measurement|243.1663773003 47.1994065115 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
2|g (SDSS PSF) AB     | 17.325    |+/-0.023|asinh mag           |6.17E+14|  4.27E-04|+/-9.04E-06|Jy|2007SDSS6.C...0000:|based on count statistics only|4858       A         | Broad-band measurement|243.1663773003 47.1994065115 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; INTERP - object contains interpolated-over pixels; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding; INTERP_CENTER - interpolated pixel(s) within 3 pixels of center; PSF_FLUX_INTERP - a signifcant amount of PSF's flux is interpolated;|From new raw data
3|r (SDSS PSF) AB     | 17.282    |+/-0.011|asinh mag           |4.77E+14|  4.44E-04|+/-4.50E-06|Jy|2007SDSS6.C...0000:|based on count statistics only|6290       A         | Broad-band measurement|243.1663773003 47.1994065115 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding; CANONICAL_BAND - this band was primary (usually r);|From new raw data
4|H{alpha} (TNG)      | 7.4E-15   |+/-20  %|erg/s/cm^2^         |4.57E+14|  7.40E+08|+/-1.48E+08|Jy-Hz|2011A&A...531A.128O|uncertainty|      6563 A         | Line measurement; flux integrated over line; lines measured in emission|16 12 39 +47 11 58 (J2000)| From fitting to map|Intermediate component flux             |From new raw data
5|H{alpha} (TNG)      | 2.0E-14   |+/-20  %|erg/s/cm^2^         |4.57E+14|  2.00E+09|+/-4.00E+08|Jy-Hz|2011A&A...531A.128O|uncertainty|      6563 A         | Line measurement; flux integrated over line; lines measured in emission|16 12 39 +47 11 58 (J2000)| From fitting to map|Broad component flux                    |From new raw data
6|i (SDSS PSF) AB     | 17.324    |+/-0.015|asinh mag           |3.89E+14|  4.27E-04|+/-5.90E-06|Jy|2007SDSS6.C...0000:|based on count statistics only|7706       A         | Broad-band measurement|243.1663773003 47.1994065115 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
7|z (SDSS PSF) AB     | 17.179    |+/-0.018|asinh mag           |3.25E+14|  4.79E-04|+/-7.94E-06|Jy|2007SDSS6.C...0000:|based on count statistics only|9222       A         | Broad-band measurement|243.1663773003 47.1994065115 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; ELLIPFAINT - no isophotal fits performed; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
8|250 GHz (IRAM/MAMBO)| 4.6E-03   |+/-0.7E-03|Jy                  |2.50E+11|  4.60E-03|+/-7.00E-04|Jy|2006AJ....132.1307P|1 sigma|     250   GHz       | Broad-band measurement|16 12 39.90 +47 11 58.0 (J2000)| Flux integrated from map|From 2003A&A...398..857O                |Averaged from previously published data; OBJ_NAME modifiedfrom published value
8|115 GHz             |           |<0.57E-03|Jy                  |2.50E+11|  |0.57E-03|Jy|2006AJ....132.1307P|1 sigma|     250   GHz       | Broad-band measurement|16 12 39.90 +47 11 58.0 (J2000)| Flux integrated from map|From 2003A&A...398..857O                |Averaged from previously published data; OBJ_NAME modifiedfrom published value
9|5.0 GHz (VLA)       ||<120E-06   |Jy                  |5.00E+09||1.20E-04|Jy|2006AJ....132.1307P|3 sigma|     5.0   GHz       | Broad-band measurement|16 12 39.90 +47 11 58.0 (J2000)| Flux integrated from map|                                        |From new raw data; OBJ_NAME modified from published value
10|1.4 GHz (VLA)       | 200E-06   |+/-20E-06|Jy                  |1.40E+09|  2.00E-04|+/-2.00E-05|Jy|2006AJ....132.1307P|1 sigma|     1.4   GHz       | Broad-band measurement|16 12 39.90 +47 11 58.0 (J2000)| Flux integrated from map|                                        |From new raw data; OBJ_NAME modified from published value
