

Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2010-09-03T10:19:38PDT



Photometric Data for SMM J163554.2+661225

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
20|450 microns (SCUBA) | 22.9      |+/-6.9 | milliJy            |6.66E+11|  22.9E-03|+/-6.9E-03|Jy|2008MNRAS.384.1611K|rms uncertainty|       450 microns   | Broad-band measurement|163554.2 +661225 (J2000)| Flux integrated from map|S/N = 12.4                              |From new raw data
20|450 microns (SCUBA) | 32        |+/-6   | milliJy            |6.66E+11|  32.0E-03|+/-6.0E-03|Jy|2008MNRAS.384.1611K|rms uncertainty|       450 microns   | Broad-band measurement|163554.2 +661225 (J2000)| Flux integrated from map|S/N = 12.4                              |From new raw data
25|850 microns (SCUBA) | 8.4       |+/-0.8 |milliJy             |3.53E+11|  8.4E-03|+/-0.8E-03|Jy|2006MNRAS.368..487K|uncertainty|     850   microns   | Broad-band measurement|163554.2 +661225 (J2000)| Flux integrated from map|                                        |From new raw data
25|850 microns (SCUBA) | 9         |+/-1   |milliJy             |3.53E+11|  9.0E-03|+/-1.0E-03|Jy|2006MNRAS.368..487K|uncertainty|     850   microns   | Broad-band measurement|163554.2 +661225 (J2000)| Flux integrated from map|                                        |From new raw data
