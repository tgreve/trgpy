
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-07-10T09:28:14PDT



Photometric Data for PKS 0156-252

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|H{alpha} (VLT)      | 1.75E-14  ||erg/s/cm^2^         |4.57E+14|  1.75E+09||Jy-Hz|2011A&A...525A..43N|no uncertainty reported|      6563 A         | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|Broad line                              |From new raw data
2|3.6 microns (IRAC)  | 291.0     |+/-29.0 | microJy            |8.44E+13|  2.91E-04|+/-2.90E-05|Jy|2007ApJS..171..353S|uncertainty|   3.550   microns   | Broad-band measurement|01 58 33.6 -24 59 31.10 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
3|4.5 microns (IRAC)  | 405.0     |+/-41.0 | microJy            |6.67E+13|  4.05E-04|+/-4.10E-05|Jy|2007ApJS..171..353S|uncertainty|   4.493   microns   | Broad-band measurement|01 58 33.6 -24 59 31.10 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
4|5.8 microns (IRAC)  | 717.0     |+/-72.0 | microJy            |5.23E+13|  7.17E-04|+/-7.20E-05|Jy|2007ApJS..171..353S|uncertainty|   5.731   microns   | Broad-band measurement|01 58 33.6 -24 59 31.10 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
5|8.0 microns (IRAC)  | 1125.0    |+/-113.0| microJy            |3.81E+13|  1.12E-03|+/-1.13E-04|Jy|2007ApJS..171..353S|uncertainty|   7.872   microns   | Broad-band measurement|01 58 33.6 -24 59 31.10 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
6|16 microns (IRS)    | 1430.0    |+/-116.6| microJy            |1.87E+13|  1.43E-03|+/-1.17E-04|Jy|2007ApJS..171..353S|uncertainty|      16   microns   | Broad-band measurement|01 58 33.6 -24 59 31.10 (J2000)| Flux in fixed aperture|6" diameter aperture                    |From reprocessed raw data
7|4.85 GHz            | 131       |+/-13   |milliJy             |4.85E+09|  1.31E-01|+/-1.30E-02|Jy|1994ApJS...90..179G|rms noise|4.85       GHz       | Broad-band measurement|015832.4 -245908 (J2000)| Modelled datum|                                        |From new raw data; Corrected for contaminating sources
8|2700 MHz            | 0.230     ||Jy                  |2.70E+09|  2.30E-01||Jy|1990PKS90.C...0000W|no uncertainty reported|    2700   MHz       | Broad-band measurement|01 56 14.0 -25 13 23 (B1950)| Integrated from scans|                                        |Homogenized from new and previously published data
9|1.4GHz              | 415.9     |+/-12.5 |milliJy             |1.40E+09|  4.16E-01|+/-1.25E-02|Jy|1998AJ....115.1693C|uncertainty|    1.40   GHz       | Broad-band measurement|01 58 33.63 -24 59 31.1 (J2000)| Flux integrated from map|High peak                               |From new raw data
10|408 MHz             | 1.39      |+/-0.05 |Jy                  |4.08E+08|  1.39E+00|+/-5.00E-02|Jy|1981MNRAS.194..693L|rms noise|408        MHz       | Broad-band measurement|015615.2 -251405 (B1950)| Modelled datum|                                        |From new raw data; Corrected for contaminating sources
11|408 MHz             | 1.390     ||Jy                  |4.08E+08|  1.39E+00||Jy|1990PKS90.C...0000W|no uncertainty reported|     408   MHz       | Broad-band measurement|01 56 14.0 -25 13 23 (B1950)| Integrated from scans|                                        |Homogenized from new and previously published data
12|365 MHz (Texas)     | 1.450     |+/-0.046|Jy                  |3.65E+08|  1.45E+00|+/-4.60E-02|Jy|1996AJ....111.1945D|internal error|365        MHz       | Broad-band measurement; obtained by interpolation over frequency|015615.163 -251405.00 (B1950)| Integrated from scans|Model:P;MFlag:C;EFlag:+;LFlag:+.        |From new raw data
13|74 MHz (VLA)        | 6.17      |+/-0.65 | Jy                 |7.38E+07|  6.17E+00|+/-6.50E-01|Jy|2007AJ....134.1245C|rms uncertainty|    73.8   MHz       | Broad-band measurement|01 58 33.33 -24 59 36.3 (J2000)| Flux integrated from map|Corrected for clean bias                |From new raw data
