
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-07-10T03:57:34PDT



Photometric Data for SDSS J100038.01+020822.4

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
2|2-10 keV (XMM)      | 8.22E-15  |+/-1.40E-15| erg/cm^2^/s        |1.45E+18|  5.67E-10|+/-9.66E-11|Jy|2007ApJS..172...29H|rms uncertainty|      6.00 keV       | Broad-band measurement|150.15809 +02.13941 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
3|2-10 keV (XMM)      | 1.02E-14  |+/-0.18E-14| erg/cm^2^/s        |1.45E+18|  7.03E-10|+/-1.24E-10|Jy|2009A&A...497..635C|statistical error|      6.00 keV       | Broad-band measurement|150.158061 +02.139463 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
4|2-10 keV (Chandra)  | 8.1E-15   |+/-1.3E-15|erg/cm^2^/s         |1.45E+18|  5.59E-10|+/-8.97E-11|Jy|2009ApJS..184..158E|uncertainty|      6.00 keV       | Broad-band measurement|150.15832 +02.13953 (J2000)| Modelled datum|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
5|0.5-10 keV (Chandra)| 1.4E-14   |+/-1.1E-15|erg/cm^2^/s         |1.27E+18|  1.10E-09|+/-8.66E-11|Jy|2009ApJS..184..158E|uncertainty|      5.25 keV       | Broad-band measurement|150.15832 +02.13953 (J2000)| Modelled datum|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
6|0.5-2 keV (XMM)     | 2.59E-15  |+/-3.07E-16| erg/cm^2^/s        |3.02E+17|  8.58E-10|+/-1.02E-10|Jy|2007ApJS..172...29H|rms uncertainty|      1.25 keV       | Broad-band measurement|150.15809 +02.13941 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
7|0.5-2 keV (XMM)     | 0.24E-14  |+/-0.02E-14| erg/cm^2^/s        |3.02E+17|  7.95E-10|+/-6.62E-11|Jy|2009A&A...497..635C|statistical error|      1.25 keV       | Broad-band measurement|150.158061 +02.139463 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
8|0.5-2 keV (Chandra) | 4.0E-15   |+/-3.6E-16|erg/cm^2^/s         |3.02E+17|  1.32E-09|+/-1.19E-10|Jy|2009ApJS..184..158E|uncertainty|      1.25 keV       | Broad-band measurement|150.15832 +02.13953 (J2000)| Modelled datum|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
9|u (SDSS PSF) AB     | 21.259    |+/-0.116|asinh mag           |8.36E+14|  1.18E-05|+/-1.26E-06|Jy|2007SDSS6.C...0000:|based on count statistics only|3585       A         | Broad-band measurement|150.1583860884 2.1395570467 (J2000)| Modelled datum|SDSS flags: MANYPETRO - more than one Petrosian radius; BAD_RADIAL - some low S/N radial points; PETROFAINT - Petrosian radius measured at very low surface brightness; ELLIPFAINT - no isophotal fits performed; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
10|g (SDSS PSF) AB     | 20.953    |+/-0.040|asinh mag           |6.17E+14|  1.51E-05|+/-5.56E-07|Jy|2007SDSS6.C...0000:|based on count statistics only|4858       A         | Broad-band measurement|150.1583860884 2.1395570467 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
11|r (SDSS PSF) AB     | 20.728    |+/-0.039|asinh mag           |4.77E+14|  1.86E-05|+/-6.67E-07|Jy|2007SDSS6.C...0000:|based on count statistics only|6290       A         | Broad-band measurement|150.1583860884 2.1395570467 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding; CANONICAL_BAND - this band was primary (usually r);|From new raw data
12|i (SDSS PSF) AB     | 20.453    |+/-0.045|asinh mag           |3.89E+14|  2.39E-05|+/-9.92E-07|Jy|2007SDSS6.C...0000:|based on count statistics only|7706       A         | Broad-band measurement|150.1583860884 2.1395570467 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
13|i (CFHT) AB         | 20.32     ||mag                 |3.86E+14|  2.70E-05||Jy|2009ApJ...696.1195T|no uncertainty reported|      7776 A         | Broad-band measurement|150.15836 +02.13961 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
14|I (HST) AB          | 20.45     ||mag                 |3.69E+14|  2.40E-05||Jy|2010ApJ...708..137M|no uncertainty reported|      8117 A         | Broad-band measurement|150.158371 +02.139555 (J2000)| Not reported in paper|                                        |Averaged from previously published data
15|F814W (HST) AB      | 20.45     || mag                |3.60E+14|  2.40E-05||Jy|2009ApJS..184..218L|no uncertainty reported|      8333 A         | Broad-band measurement|150.158371 +02.139555 (J2000)| Total flux|                                        |From new raw data
16|F814W (HST/ACS) AB      | 20.21     || mag                |3.60E+14|  2.99E-05||Jy|2007ApJS..172..383T|no uncertainty reported|      8333 A         | Broad-band measurement|150.1583557 +02.1396151 (J2000)| Not reported in paper|S/N = 15.81                             |Averaged from previously published data
17|z (SDSS PSF) AB     | 20.366    |+/-0.194|asinh mag           |3.25E+14|  2.52E-05|+/-4.60E-06|Jy|2007SDSS6.C...0000:|based on count statistics only|9222       A         | Broad-band measurement|150.1583860884 2.1395570467 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; ELLIPFAINT - no isophotal fits performed; BINNED1 - detected at >=5 sigma in original imaging frame;|From new raw data
18|3.6 microns (IRAC)  | 116.915   |+/-0.180| microJy            |8.44E+13|  1.17E-04|+/-1.80E-07|Jy|2009AJ....137.3884R|uncertainty|     3.550 microns   | Broad-band measurement|150.158386 2.139557 (J2000)| Flux integrated from map|                                        |From new raw data
19|4.5 microns (IRAC)  | 174.770   |+/-0.280| microJy            |6.67E+13|  1.75E-04|+/-2.80E-07|Jy|2009AJ....137.3884R|uncertainty|     4.493 microns   | Broad-band measurement|150.158386 2.139557 (J2000)| Flux integrated from map|                                        |From new raw data
20|5.8 microns (IRAC)  | 257.968   |+/-0.750| microJy            |5.23E+13|  2.58E-04|+/-7.50E-07|Jy|2009AJ....137.3884R|uncertainty|     5.731 microns   | Broad-band measurement|150.158386 2.139557 (J2000)| Flux integrated from map|                                        |From new raw data
21|8.0 microns (IRAC)  | 354.672   |+/-1.360| microJy            |3.81E+13|  3.55E-04|+/-1.36E-06|Jy|2009AJ....137.3884R|uncertainty|     7.872 microns   | Broad-band measurement|150.158386 2.139557 (J2000)| Flux integrated from map|                                        |From new raw data
22|24 microns (MIPS)   | 1.59      ||milliJy             |1.27E+13|  1.59E-03||Jy|2010ApJ...716..348B|no uncertainty reported|     23.68 microns   | Broad-band measurement|150.1583900 2.1396030 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
23|[C II] 158 (CSO)    | 1.74E-18  |+/-0.40E-18|W/m^2^              |1.90E+12|  1.74E+08|+/-4.00E+07|Jy-Hz|2010ApJ...724..957S|statistical error|       158 microns   | Line measurement; flux integrated over line; lines measured in emission|10 00 38.0 +02 08 22.4 (J2000)| Flux integrated from map|                                        |From new raw data
24|244.603 GHz (IRAM)  | 10.35     ||milliJy             |2.45E+11|  1.03E-02||Jy|2008A&A...491..173A|no uncertainty reported|   244.603 GHz       | Broad-band measurement|10 00 38.01 +02 08 22.6 (J2000)| Flux integrated from map|                                        |From new raw data
25|203.850 GHz (IRAM)  | 11.56     ||milliJy             |2.04E+11|  1.16E-02||Jy|2008A&A...491..173A|no uncertainty reported|   203.850 GHz       | Broad-band measurement|10 00 38.01 +02 08 22.6 (J2000)| Flux integrated from map|                                        |From new raw data
26|163.088 GHz (IRAM)  | 8.39      ||milliJy             |1.63E+11|  8.39E-03||Jy|2008A&A...491..173A|no uncertainty reported|   163.088 GHz       | Broad-band measurement|10 00 38.01 +02 08 22.6 (J2000)| Flux integrated from map|                                        |From new raw data
27|81.551 GHz (IRAM)   | 3.08      ||milliJy             |8.16E+10|  3.08E-03||Jy|2008A&A...491..173A|no uncertainty reported|    81.551 GHz       | Broad-band measurement|10 00 38.01 +02 08 22.6 (J2000)| Flux integrated from map|                                        |From new raw data
28|1.4 GHz (VLA)       | 237       |+/-27   | microJy            |1.40E+09|  2.37E-04|+/-2.70E-05|Jy|2007ApJS..172..132B|uncertainty|      1.40 GHz       | Broad-band measurement|10 00 38.02 +02 08 22.6 (J2000)| Flux integrated from map|                                        |From new raw data
29|1.4 GHz (VLA)       | 0.237     |+/-0.027| milliJy            |1.40E+09|  2.37E-04|+/-2.70E-05|Jy|2007ApJS..172...46S|statistical error|       1.4 GHz       | Broad-band measurement|10 00 38.016 +02 08 22.56 (J2000)| Flux integrated from map|                                        |From new raw data
30|1.4 GHz (VLA)       | 0.272     |+/-0.083|milliJy             |1.40E+09|  2.72E-04|+/-8.30E-05|Jy|2004AJ....128.1974S|uncertainty|     1.4   GHz       | Broad-band measurement|10 00 38.022 +02 08 22.85 (J2000)| Flux integrated from map|                                        |From new raw data
31|1.4 GHz (VLA)       | 175       |+/-8    | microJy            |1.40E+09|  1.75E-04|+/-8.00E-06|Jy|2007ApJS..172..132B|uncertainty|      1.40 GHz       | Broad-band measurement|10 00 38.02 +02 08 22.6 (J2000)| Peak flux|                                        |From new raw data
