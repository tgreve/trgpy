
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-06-17T16:37:41PDT



Photometric Data for BzK 04171

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|3.6 microns (IRAC)  | 24.00     |+/-1.20 |microJy             |8.44E+13|  2.40E-05|+/-1.20E-06|Jy|2011AJ....141....1T|rms uncertainty|     3.550 microns   | Broad-band measurement|189.110626 62.143169 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
2|4.5 microns (IRAC)  | 27.90     |+/-1.40 |microJy             |6.67E+13|  2.79E-05|+/-1.40E-06|Jy|2011AJ....141....1T|rms uncertainty|     4.493 microns   | Broad-band measurement|189.110626 62.143169 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
3|5.8 microns (IRAC)  | 23.10     |+/-1.24 |microJy             |5.23E+13|  2.31E-05|+/-1.24E-06|Jy|2011AJ....141....1T|rms uncertainty|     5.731 microns   | Broad-band measurement|189.110626 62.143169 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
4|8.0 microns (IRAC)  | 22.00     |+/-1.23 |microJy             |3.81E+13|  2.20E-05|+/-1.23E-06|Jy|2011AJ....141....1T|rms uncertainty|     7.872 microns   | Broad-band measurement|189.110626 62.143169 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
5|16 microns (IRS)    | 125.2     |+/-15.0 |microJy             |1.90E+13|  1.25E-04|+/-1.50E-05|Jy|2011AJ....141....1T|rms uncertainty|      15.8 microns   | Broad-band measurement|189.110626 62.143169 (J2000)| From fitting to map|                                        |From new raw data
6|24 microns (MIPS)   | 139.0     |+/-6.4  |microJy             |1.27E+13|  1.39E-04|+/-6.40E-06|Jy|2011AJ....141....1T|rms uncertainty|     23.68 microns   | Broad-band measurement|189.110626 62.143169 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
7|24 microns (MIPS)   | 142       ||microJy             |1.27E+13|  1.42E-04||Jy|2011ApJ...726...93R|no uncertainty reported|     23.68 microns   | Broad-band measurement|12 36 26.52 +62 08 35.4 (J2000)| Not reported in paper|                                        |Averaged from previously published data
8|24 microns (MIPS)   | 148.5     |+/-5.6  |microJy             |1.27E+13|  1.49E-04|+/-5.60E-06|Jy|2011A&A...528A..35M|uncertainty|     23.68 microns   | Broad-band measurement|12 36 26.55 +62 08 35.34 (J2000)| Flux integrated from map|                                        |From new raw data
9|70 microns (MIPS)   ||<5.8       |milliJy             |4.20E+12||5.80E-03|Jy|2011A&A...528A..35M|no uncertainty reported|     71.42 microns   | Broad-band measurement|12 36 26.55 +62 08 35.34 (J2000)| Flux integrated from map|                                        |From new raw data
10|CO(3-2) (IRAM)      | 0.70      |+/-0.15 |Jy km/s             |3.46E+11|  3.20E+05|+/-6.86E+04|Jy-Hz|2009ApJ...698L.178D|uncertainty|   345.796 GHz       | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|                                        |From new raw data
11|CO[2-1] (IRAM)      | 0.65      ||Jy km/s             |2.31E+11|  2.03E+05||Jy-Hz|2010ApJ...713..686D|no uncertainty reported|   230.538 GHz       | Line measurement; flux integrated over line; lines measured in emission|12 36 26.516 +62 08 35.35 (J2000)| Flux integrated from map|                                        |From new raw data
12|CO(2-1) (IRAM)      | 0.60      |+/-0.09 | Jy km/s            |2.31E+11|  1.87E+05|+/-2.81E+04|Jy-Hz|2008ApJ...673L..21D|uncertainty|   230.539 GHz       | Line measurement; flux integrated over line; lines measured in emission|12 36 26.53 +62 08 35.3 (J2000)| Flux integrated from map|                                        |From new raw data
13|CO(2-1) (IRAM)      | 0.62      |+/-0.07 |Jy km/s             |2.30E+11|  1.89E+05|+/-2.13E+04|Jy-Hz|2009ApJ...698L.178D|uncertainty|   230.538 GHz       | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|                                        |From new raw data
14|CO(1-0) (VLA)       | 0.20      |+/-0.05 |Jy km/s             |1.15E+11|  3.12E+04|+/-7.80E+03|Jy-Hz|2010ApJ...718..177A|uncertainty|   115.271 GHz       | Line measurement; flux integrated over line; lines measured in emission|12 36 26.516 +62 08 35.35 (J2000)| Flux integrated from map|                                        |From new raw data
15|1.4 GHz (VLA)       | 41        |+/-7    | microJy            |1.40E+09|  4.10E-05|+/-7.00E-06|Jy|2006MNRAS.371..963B|1 sigma|       1.4 GHz       | Broad-band measurement|12 36 26.547 +62 08 35.39 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
16|1.4 GHz (VLA)       | 31.3      |+/-8.1  |microJy             |1.40E+09|  3.13E-05|+/-8.10E-06|Jy|2010ApJS..188..178M|uncertainty|       1.4 GHz       | Broad-band measurement|12 36 26.52 +62 08 35.3 (J2000)| Total flux; Beam filling or dilution corrected|Major=0.9"; Minor=0.0"; PA=178 deg      |From new raw data
