
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-04-05T08:15:36PDT



Photometric Data for SMMJ021738-050339

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|850 microns (SCUBA) | 4.4       |+/-1.7  | milliJy            |3.53E+11|4.4E-03|+/-1.7E-03|Jy|2004ApJ...614..671C|1 sigma|       850 microns   | Broad-band measurement|163656.28 +405912.2 (J2000)| Flux integrated from map|                                        |From new raw data
2|1.4 GHz (VLA)       | 57       |+/-10   | microJy            |1.40E+09|  57.E-06|+/-10.E-06|Jy|2006MNRAS.371..963B|1 sigma|       1.4 GHz       | Broad-band measurement|16 36 55.767 +40 59 09.97 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
