


Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.





Photometric Data 

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|4.5um (Spitzer) | 10.1  |+/-1.0| uJy  | 6.67E13| 10.1E-6| 1.0E-6 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
2|8.0um (Spitzer) | 15.4 |+/-1.5| uJy  | 3.75E13| 15.4E-6| 1.5E-6 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
3|24um (Spitzer)  | 12.0 |+/-4.3| uJy  | 1.25E13| 12.0E-6| 4.3E-6 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
4|850um (SCUBA)   | 9.9 |+/-2.3| mJy  | 3.529E11| 9.9E-3| 2.3E-3 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
5|2mm (PdBI)      | 0.20|+/-0.06|mJy  | 136.96E9| 0.30E-03|+/-0.1E-03 |Jy |2003MNRAS.343..293M|rms uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
6|3.3mm (PdBI)    |  |<0.18| mJy  | 9.09E10| |0.18E-03 |Jy |2003MNRAS.343..293M|3rms uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
7|1.4GHz (VLA)    | 32.2 |+/-6.5| uJy  | 1.4E9| 32.3E-6| 6.5E-6 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
