
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-06-17T16:58:46PDT



Photometric Data for PKS 0114-21

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|3.6 microns (IRAC)  | 87.3      |+/-8.9  | microJy            |8.44E+13|  8.73E-05|+/-8.90E-06|Jy|2007ApJS..171..353S|uncertainty|   3.550   microns   | Broad-band measurement|01 16 51.4 -20 52 06.71 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
2|4.5 microns (IRAC)  | 117.0     |+/-12.0 | microJy            |6.67E+13|  1.17E-04|+/-1.20E-05|Jy|2007ApJS..171..353S|uncertainty|   4.493   microns   | Broad-band measurement|01 16 51.4 -20 52 06.71 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
3|5.8 microns (IRAC)  | 157.0     |+/-16.0 | microJy            |5.23E+13|  1.57E-04|+/-1.60E-05|Jy|2007ApJS..171..353S|uncertainty|   5.731   microns   | Broad-band measurement|01 16 51.4 -20 52 06.71 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
4|8.0 microns (IRAC)  | 398.0     |+/-40.0 | microJy            |3.81E+13|  3.98E-04|+/-4.00E-05|Jy|2007ApJS..171..353S|uncertainty|   7.872   microns   | Broad-band measurement|01 16 51.4 -20 52 06.71 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
5|22 GHz (ATCA)       | 0.243     |+/-0.024|Jy                  |2.20E+10|  2.43E-01|+/-2.40E-02|Jy|2006A&A...445..465R|uncertainty|      22   GHz       | Broad-band measurement|| Modelled datum|                                        |From new raw data
6|20 GHz (ATCA)       | 240       |+/-16   |milliJy             |1.99E+10|  2.40E-01|+/-1.60E-02|Jy|2010MNRAS.402.2403M|rms uncertainty|    19.904 GHz       | Broad-band measurement|01 16 51.47 -20 52 06.5 (J2000)| Flux integrated from map|                                        |From new raw data
7|18.5 GHz (ATCA)     | 0.283     |+/-0.014|Jy                  |1.85E+10|  2.83E-01|+/-1.40E-02|Jy|2006A&A...445..465R|uncertainty|    18.5   GHz       | Broad-band measurement|| Modelled datum|                                        |From new raw data
8|10695 MHz           | 0.54      |+/-.01  |Jy                  |1.07E+10|  5.40E-01|+/-1.00E-02|Jy|1981A&AS...45..367K|uncertainty|   10695   MHz       | Broad-band measurement|011425.91 -210753.4 (B1950)| Not reported in paper|                                        |From new raw data
9|8870 MHz            | 0.66      |+/-.03  |Jy                  |8.87E+09|  6.60E-01|+/-3.00E-02|Jy|1973AuJPh..26...93S|uncertainty|    8870   MHz       | Broad-band measurement|011425.91 -210753.4 (B1950)| Not reported in paper|From Kuhr catalog (1981A&AS...45..367K) |Transformed from previously published data
10|8400 MHz            | 0.67      ||Jy                  |8.40E+09|  6.70E-01||Jy|1990PKS90.C...0000W|no uncertainty reported|    8400   MHz       | Broad-band measurement|01 14 26.0 -21 07 55 (B1950)| Integrated from scans|                                        |Homogenized from new and previously published data
11|8 GHz (ATCA)        | 750       |+/-39   |milliJy             |8.00E+09|  7.50E-01|+/-3.90E-02|Jy|2010MNRAS.402.2403M|rms uncertainty|         8 GHz       | Broad-band measurement|01 16 51.47 -20 52 06.5 (J2000)| Flux integrated from map|                                        |From new raw data
12|5009 MHz            | 1.28      |+/-.08  |Jy                  |5.01E+09|  1.28E+00|+/-8.00E-02|Jy|1981A&AS...45..367K|uncertainty|    5009   MHz       | Broad-band measurement|011425.91 -210753.4 (B1950)| Not reported in paper|Recal. to Baars scale by factor of 1.03 |Recalibrated data
13|5000 MHz            | 1.240     ||Jy                  |5.00E+09|  1.24E+00||Jy|1990PKS90.C...0000W|no uncertainty reported|    5000   MHz       | Broad-band measurement|01 14 26.0 -21 07 55 (B1950)| Integrated from scans|                                        |Homogenized from new and previously published data
14|5 GHz (ATCA)        | 1661      |+/-83   |milliJy             |5.00E+09|  1.66E+00|+/-8.30E-02|Jy|2010MNRAS.402.2403M|rms uncertainty|         5 GHz       | Broad-band measurement|01 16 51.47 -20 52 06.5 (J2000)| Flux integrated from map|                                        |From new raw data
15|4.85 GHz            | 1415      |+/-74   |milliJy             |4.85E+09|  1.42E+00|+/-7.40E-02|Jy|1994ApJS...90..179G|rms noise|4.85       GHz       | Broad-band measurement|011650.9 -205210 (J2000)| Modelled datum|                                        |From new raw data; Corrected for contaminating sources
16|2700 MHz            | 2.23      |+/-.09  |Jy                  |2.70E+09|  2.23E+00|+/-9.00E-02|Jy|1976AuJPA..39....1W|uncertainty|    2700   MHz       | Broad-band measurement|011425.91 -210753.4 (B1950)| Not reported in paper|From Kuhr catalog (1981A&AS...45..367K) |Transformed from previously published data
17|2700 MHz            | 2.400     ||Jy                  |2.70E+09|  2.40E+00||Jy|1990PKS90.C...0000W|no uncertainty reported|    2700   MHz       | Broad-band measurement|01 14 26.0 -21 07 55 (B1950)| Integrated from scans|                                        |Homogenized from new and previously published data
18|2650 MHz            | 2.22      |+/-.05  |Jy                  |2.65E+09|  2.22E+00|+/-5.00E-02|Jy|1975AuJPA..38....1W|uncertainty|    2650   MHz       | Broad-band measurement|011425.91 -210753.4 (B1950)| Not reported in paper|From Kuhr catalog (1981A&AS...45..367K) |Transformed from previously published data
19|1410 MHz            | 4.100     ||Jy                  |1.41E+09|  4.10E+00||Jy|1990PKS90.C...0000W|no uncertainty reported|    1410   MHz       | Broad-band measurement|01 14 26.0 -21 07 55 (B1950)| Integrated from scans|                                        |Homogenized from new and previously published data
20|1410 MHz            | 4.22      |+/-.06  |Jy                  |1.41E+09|  4.22E+00|+/-6.00E-02|Jy|1981A&AS...45..367K|uncertainty|    1410   MHz       | Broad-band measurement|011425.91 -210753.4 (B1950)| Not reported in paper|Recal. to Baars scale by factor of 1.017|Recalibrated data
21|1.4GHz              | 4091.6    |+/-122.7|milliJy             |1.40E+09|  4.09E+00|+/-1.23E-01|Jy|1998AJ....115.1693C|uncertainty|    1.40   GHz       | Broad-band measurement|01 16 51.43 -20 52 6.6 (J2000)| Flux integrated from map|                                        |From new raw data
22|960 MHz             | 5.75      |+/-.11  |Jy                  |9.60E+08|  5.75E+00|+/-1.10E-01|Jy|1981A&AS...45..367K|uncertainty|     960   MHz       | Broad-band measurement|011425.91 -210753.4 (B1950)| Not reported in paper|Recal. to Baars scale by factor of 1.029|Recalibrated data
23|635 MHz             | 8.04      |+/-.21  |Jy                  |6.35E+08|  8.04E+00|+/-2.10E-01|Jy|1981A&AS...45..367K|uncertainty|     635   MHz       | Broad-band measurement|011425.91 -210753.4 (B1950)| Not reported in paper|Recal. to Baars scale by factor of 1.035|Recalibrated data
24|468 MHz             | 10.2      |+/-.26  |Jy                  |4.68E+08|  1.02E+01|+/-2.60E-01|Jy|1981A&AS...45..367K|uncertainty|     468   MHz       | Broad-band measurement|011425.91 -210753.4 (B1950)| Not reported in paper|Recal. to Baars scale by factor of 1.045|Recalibrated data
25|408 MHz             | 10.60     ||Jy                  |4.08E+08|  1.06E+01||Jy|1990PKS90.C...0000W|no uncertainty reported|     408   MHz       | Broad-band measurement|01 14 26.0 -21 07 55 (B1950)| Integrated from scans|                                        |Homogenized from new and previously published data
26|408 MHz             | 10.64     |+/-0.23 |Jy                  |4.08E+08|  1.06E+01|+/-2.30E-01|Jy|1981MNRAS.194..693L|rms noise|408        MHz       | Broad-band measurement|011425.9 -210754 (B1950)| Modelled datum|                                        |From new raw data; Corrected for contaminating sources
27|365 MHz             | 10.67     |+/-.63  |Jy                  |3.65E+08|  1.07E+01|+/-6.30E-01|Jy|1981A&AS...45..367K|uncertainty|     365   MHz       | Broad-band measurement|011425.91 -210753.4 (B1950)| Not reported in paper|Recal. to Baars scale by factor of 1.047|Recalibrated data
28|365 MHz (Texas)     | 11.033    |+/-0.179|Jy                  |3.65E+08|  1.10E+01|+/-1.79E-01|Jy|1996AJ....111.1945D|internal error|365        MHz       | Broad-band measurement; obtained by interpolation over frequency|011426.011 -210754.77 (B1950)| Integrated from scans|Model:P;MFlag:+;EFlag:+;LFlag:+.        |From new raw data
29|160 MHz             | 15.3      ||Jy                  |1.60E+08|  1.53E+01||Jy|1995AuJPh..48..143S|no uncertainty reported|160        MHz       | Broad-band measurement|011424.6 -210753. (B1950)| Flux integrated from map|                                        |From new raw data
30|145 MHz (PAPER)     | 12.0      ||Jy                  |1.45E+08|  1.20E+01||Jy|2011ApJ...734L..34J|no uncertainty reported|       145 MHz       | Broad-band measurement|19.25 -20.74 (J2000)| Flux integrated from map|                                        |From new raw data
31|80 MHz              | 18.       ||Jy                  |8.00E+07|  1.80E+01||Jy|1995AuJPh..48..143S|no uncertainty reported| 80        MHz       | Broad-band measurement|011424.6 -210753. (B1950)| Flux integrated from map|                                        |From new raw data
32|80 MHz              | 18.00     ||Jy                  |8.00E+07|  1.80E+01||Jy|1990PKS90.C...0000W|no uncertainty reported|      80   MHz       | Broad-band measurement|01 14 26.0 -21 07 55 (B1950)| Integrated from scans|                                        |Homogenized from new and previously published data
33|74 MHz (VLA)        | 13.76     |+/-1.40 | Jy                 |7.38E+07|  1.38E+01|+/-1.40E+00|Jy|2007AJ....134.1245C|rms uncertainty|    73.8   MHz       | Broad-band measurement|01 16 51.40 -20 52 09.1 (J2000)| Flux integrated from map|Corrected for clean bias                |From new raw data
