
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-05-28T01:42:09PDT



Photometric Data for PEPJ123634+620627 (z=1.215)

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|R (Keck II) AB      | 24.36     || mag                |4.62E+14|  6.55E-07||Jy|2004AJ....127.3121W|no uncertainty reported|   648.7   A         | Broad-band measurement|12 36 34.531 +62 06 27.78 (J2000)| Total flux|                                        |From new raw data
2|3.6 microns (IRAC)  | 70.60     |+/-3.53 |microJy             |8.44E+13|  7.06E-05|+/-3.53E-06|Jy|2011AJ....141....1T|rms uncertainty|     3.550 microns   | Broad-band measurement|189.143692 62.107803 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
3|4.5 microns (IRAC)  | 64.70     |+/-3.24 |microJy             |6.67E+13|  6.47E-05|+/-3.24E-06|Jy|2011AJ....141....1T|rms uncertainty|     4.493 microns   | Broad-band measurement|189.143692 62.107803 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
4|5.8 microns (IRAC)  | 47.00     |+/-2.40 |microJy             |5.23E+13|  4.70E-05|+/-2.40E-06|Jy|2011AJ....141....1T|rms uncertainty|     5.731 microns   | Broad-band measurement|189.143692 62.107803 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
5|8.0 microns (IRAC)  | 39.80     |+/-2.08 |microJy             |3.81E+13|  3.98E-05|+/-2.08E-06|Jy|2011AJ....141....1T|rms uncertainty|     7.872 microns   | Broad-band measurement|189.143692 62.107803 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
6|16 microns (IRS)    | 167.0     |+/-19.8 |microJy             |1.90E+13|  1.67E-04|+/-1.98E-05|Jy|2011AJ....141....1T|rms uncertainty|      15.8 microns   | Broad-band measurement|189.143692 62.107803 (J2000)| From fitting to map|                                        |From new raw data
1|MIPS 24 microns      | 108.      |+/-9.0  |microJy         |1.25E+13   |  108.E-06|+/-9.0E-06  |Jy|1990IRASF.C...0000M|3sigma uncertainty| 25        microns   | Broad-band measurement|115813.1 +302058 (B1950)| Flux in fixed aperture|                                        |From new raw data
8|24 microns (MIPS)   | 96.3      |+/-6.2  |microJy             |1.27E+13|  9.63E-05|+/-6.20E-06|Jy|2011A&A...528A..35M|uncertainty|     23.68 microns   | Broad-band measurement|12 36 34.49 +62 06 28.02 (J2000)| Flux integrated from map|                                        |From new raw data
2|70 microns (PACS)    |           |<2.0    |mJy             |4.283e+12  |          |2.0E-03     |Jy|2.40e+01           |3sigma |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
9|70 microns (MIPS)   ||<2.8       |milliJy             |4.20E+12||2.80E-03|Jy|2011A&A...528A..35M|3sigma |     71.42 microns   | Broad-band measurement|12 36 34.49 +62 06 28.02 (J2000)| Flux integrated from map|                                        |From new raw data
3|100 microns (PACS)   | 7.1       |+/-0.4  |mJy             |2.998e+12  |  7.1E-03 |+/-0.4E-03  |Jy|2.40e+01           |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
4|160 microns (PACS)   | 13.4      |+/-1.2  |mJy             |1.874e+12  | 13.4E-03 |+/-1.2E-03  |Jy|2.40e+01           |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
5|250 microns (SPIRE)  | 18.1      |+/-4.0  |mJy             |1.199e+12  |  18.1E-03|+/-4.0e-03  |Jy|2.40e+01           |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
6|350 microns (SPIRE)  | 16.1      |+/-3.0  |mJy             |8.565e+11  |  16.1E-03|+/-3.0e-03  |Jy|2.40e+01           |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
7|500 microns (SPIRE)  | 15.1      |+/-4.0  |mJy             |5.996e+11  |  15.1E-03|+/-4.0e-03  |Jy|2.40e+01           |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
8|1160 microns (Penner)|           |<2.0    |mJy             |2.58442E+11|          |2.0E-03     |Jy|2004MNRAS.354..779G|3sigma uncertainty|      1200 microns   | Broad-band measurement|16 36 55.9 +40 59 12 (J2000)| Flux integrated from map|S/N = 3.66                              |From new raw data
10|1.4 GHz (VLA)       | 27.5      |+/-5.1  |microJy             |1.40E+09|  2.75E-05|+/-5.10E-06|Jy|2010ApJS..188..178M|uncertainty|       1.4 GHz       | Broad-band measurement|12 36 34.49 +62 06 28.1 (J2000)| Total flux; Beam filling or dilution corrected|Major=0.0"; Minor=0.0"; PA=0 deg        |From new raw data
