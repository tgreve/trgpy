
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-07-10T03:41:13PDT



Photometric Data for [HB89] 0957+561

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|F555W (HST/WFPC2)         | 19.05     |+/-0.06 | mag                |5.54E+14|  8.95E-05|+/-4.95E-06|Jy|2008A&A...478...95Y|uncertainty|      5407 A         | Broad-band measurement|| Modelled datum|                                        |Averaged from previously published data
2|F606W (HST) AB      | 18.809    |+/-0.061|mag                 |4.97E+14|  1.09E-04|+/-6.11E-06|Jy|2010ApJ...711..246F|uncertainty|      6033 A         | Broad-band measurement|| Total flux|                                        |From new raw data
3|F814W (HST/WFPC2)         | 17.12     |+/-0.03 | mag                |3.78E+14|  3.53E-04|+/-9.76E-06|Jy|2008A&A...478...95Y|uncertainty|      7940 A         | Broad-band measurement|| Modelled datum|                                        |Averaged from previously published data
4|F814W (HST/ACS) AB      | 17.743    |+/-0.065|mag                 |3.68E+14|  2.90E-04|+/-1.74E-05|Jy|2010ApJ...711..246F|uncertainty|      8140 A         | Broad-band measurement|| Total flux|                                        |From new raw data
5|I (HST)             | 15.99     ||mag                 |3.68E+14|  9.68E-04||Jy|2011ApJ...738...96M|no uncertainty reported|     0.814 microns   | Broad-band measurement|| Not reported in paper|                                        |From reprocessed raw data
6|F160W (HST/NIC2)    | 17.05     ||mag                 |1.87E+14|  1.64E-04||Jy|2006ApJ...649..616P|no uncertainty reported|   1.606   microns   | Broad-band measurement|10 01 20.78 +55 53 49.4 (J2000)| From fitting to map|Quasar mag; extinction = 0.01           |From new raw data; Extinction-corrected for Milky Way
7|F160W (HST/NIC2)    | 17.83     |+/-0.3  |mag                 |1.87E+14|  7.99E-05|+/-4.31E-06|Jy|2006ApJ...649..616P|typical accuracy|   1.606   microns   | Broad-band measurement|10 01 20.78 +55 53 49.4 (J2000)| From fitting to map|Host mag; extinction = 0.01             |From new raw data; Extinction-corrected for Milky Way
8|F160W (HST)         | 15.14     |+/-0.09 | mag                |1.87E+14|  9.17E-04|+/-7.60E-05|Jy|2008A&A...478...95Y|uncertainty|     1.603 microns   | Broad-band measurement|| Modelled datum|                                        |Averaged from previously published data
9|F160W (HST)         | 16.51     ||mag                 |1.87E+14|  2.60E-04||Jy|2011ApJ...742...93A|no uncertainty reported|      1.60 microns   | Broad-band measurement|| Not reported in paper|Unmagnified quasar mag                  |Averaged from previously published data
10|8.4 GHz (VLBI)      | 11        ||milliJy             |8.40E+09|  1.10E-02||Jy|2010A&A...520A.113B|no uncertainty reported|       8.4 GHz       | Broad-band measurement|10 01 20.6911 +55 53 55.611 (J2000)| Flux integrated from map|Correlated flux                         |From new raw data
11|5 GHz (VLA)         | 51        ||milliJy             |4.89E+09|  5.10E-02||Jy|1997A&AS..122..235L|no uncertainty reported|     4.885 GHz       | Broad-band measurement|10 01 21.32 +55 53 58.1 (J2000)| Flux integrated from map|Core flux; S/N = 57                     |From new raw data
12|4.85 GHz            | 205       |+/-22   |milliJy             |4.85E+09|  2.05E-01|+/-2.20E-02|Jy|1991ApJS...75.1011G|rms noise|4.85       GHz       | Broad-band measurement|095758.5 +560808 (B1950)| Modelled datum|                                        |From new raw data; Corrected for contaminating sources
13|4.85 GHz            | 203       |+/-15  %|milliJy             |4.85E+09|  2.03E-01|+/-3.05E-02|Jy|1991ApJS...75....1B|uncertainty|4.85       GHz       | Broad-band measurement|095759.5 +560812 (B1950)| Peak flux|                                        |From new raw data; Corrected for contaminating sources
14|2.3 GHz (VLBI)      | 24        ||milliJy             |2.30E+09|  2.40E-02||Jy|2010A&A...520A.113B|no uncertainty reported|       2.3 GHz       | Broad-band measurement|10 01 20.6911 +55 53 55.611 (J2000)| Flux integrated from map|Correlated flux                         |From new raw data
15|1.40 GHz            | 494       ||milliJy             |1.40E+09|  4.94E-01||Jy|1992ApJS...79..331W|no uncertainty reported|1.4        GHz       | Broad-band measurement|095759.5 +560812 (B1950)| Peak flux|                                        |From new raw data
16|1.4GHz (VLA)             | 551.9     |+/-16.6 |milliJy             |1.40E+09|  5.52E-01|+/-1.66E-02|Jy|1998AJ....115.1693C|uncertainty|    1.40   GHz       | Broad-band measurement|10 01 21.07 +55 53 55.8 (J2000)| Flux integrated from map|                                        |From new raw data
17|365 MHz (Texas)     | 1.628     |+/-0.030|Jy                  |3.65E+08|  1.63E+00|+/-3.00E-02|Jy|1996AJ....111.1945D|internal error|365        MHz       | Broad-band measurement; obtained by interpolation over frequency|095757.562 560823.50 (B1950)| Integrated from scans|Model:P;MFlag:+;EFlag:C;LFlag:+.        |From new raw data
18|151 MHz (6C)        | 2.91      |+/-0.040|Jy                  |1.52E+08|  2.91E+00|+/-4.00E-02|Jy|1990MNRAS.246..256H|typical accuracy|151.5      MHz       | Broad-band measurement|095757.6 560821. (B1950)| Peak flux|                                        |From new raw data
19|151 MHz (6C)        | 2.85      |+/-0.090|Jy                  |1.52E+08|  2.85E+00|+/-9.00E-02|Jy|1990MNRAS.246..256H|typical accuracy|151.5      MHz       | Broad-band measurement|095757.6 560821. (B1950)| Flux integrated from map|                                        |From new raw data
20|74 MHz (VLA)        | 4.37      |+/-0.44 | Jy                 |7.38E+07|  4.37E+00|+/-4.40E-01|Jy|2007AJ....134.1245C|rms uncertainty|      73.8 MHz       | Broad-band measurement|10 01 20.88 +55 53 53.9 (J2000)| Flux integrated from map|Corrected for clean bias                |From new raw data
21|38 MHz (8C)         | 7.5       |+/-15.0%|Jy                  |3.78E+07|  7.50E+00|+/-1.12E+00|Jy|1995MNRAS.274..447H|no uncertainty reported|38         MHz       | Broad-band measurement|095800. +560903. (B1950)| Peak flux|Part of multiple component source       |From new raw data
22|38 MHz (8C)         | 8.9       |+/-1.4  |Jy                  |3.78E+07|  8.90E+00|+/-1.41E+00|Jy|1995MNRAS.274..447H|2.5 times noise|38         MHz       | Broad-band measurement|095800. +560903. (B1950)| Flux integrated from map|Part of multiple component source       |From new raw data
