

Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.


queryDateTime:2009-11-03T15:32:02PST



Photometric Data for SMM J09431+4700

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|450 microns (SCUBA) | -32       |+/-140  |milliJy             |6.66E+11| -3.20E-02|+/-1.40E-01|Jy|2007MNRAS.376.1073Z|1sigma uncertainty|     450   microns   | Broad-band measurement|09 43 05.1 +47 00 10 (J2000)| Flux integrated from map|                                        |From reprocessed raw data
2|850 microns (SCUBA) | 5.1       |+/-1.5 |milliJy             |3.53E+11|  5.1E-03|+/-1.5E-03 |Jy|2007MNRAS.376.1073Z|no uncertainty reported|     850   microns   | Broad-band measurement|09 43 05.1 +47 00 10 (J2000)| Flux integrated from map|S/N = 4.5                               |From reprocessed raw data
3|1.3 mm (PdBI)       | 2.2       |+/-0.3  |milliJy             |2.31E+11|  2.20E-03|+/-3.00E-04|Jy|2006ApJ...640..228T|uncertainty|     1.3   mm        | Broad-band measurement| | Flux integrated from map|                                        |From new raw data
4|1.1 cm (EVLA)       |        |<44.0  |microJy             |2.73E+10|  |44.E-06|Jy|2006ApJ...640..228T|3sigma uncertainty|     1.1   cm        | Broad-band measurement| | Flux integrated from map|                                        |From new raw data
5|1.4GHz  | 55.      | 10.|milliJy             |1.4E+9|  55.E-06|10.E-6 |Jy|2007MNRAS.376.1073Z|no uncertainty reported|     850   microns   | Broad-band measurement|14 01 04.7 +02 52 28 (J2000)| Flux integrated from map|S/N = 9.6                               |From reprocessed raw data
