
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-06-16T05:01:41PDT



Photometric Data for DEEP2 12004280

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|K_s (Keck)          | 18.32     || mag                |1.39E+14|  2.91E-05||Jy|2007MNRAS.382..109T|no uncertainty reported|      2.15 microns   | Broad-band measurement|214.25360 +52.45039 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
