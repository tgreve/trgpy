
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-06-16T05:48:13PDT



Photometric Data for DEEP2 13004661

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|CO(3-2) (PdBI)      ||<0.06      |Jy km/s             |3.46E+11|  1.69E+05|3.16E+04|Jy-Hz|2010Natur.463..781T|3 sigma|   345.998 GHz       | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|                                        |From new raw data
