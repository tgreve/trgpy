
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-07-10T12:48:07PDT



Photometric Data for LEDA 2823709

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|3.6 microns (IRAC)  | 23.6      |+/-2.6  | microJy            |8.44E+13|  2.36E-05|+/-2.60E-06|Jy|2007ApJS..171..353S|uncertainty|   3.550   microns   | Broad-band measurement|03 52 51.6 -27 49 22.61 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
2|4.5 microns (IRAC)  | 40.6      |+/-4.2  | microJy            |6.67E+13|  4.06E-05|+/-4.20E-06|Jy|2007ApJS..171..353S|uncertainty|   4.493   microns   | Broad-band measurement|03 52 51.6 -27 49 22.61 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
3|5.8 microns (IRAC)  | 82.2      |+/-27.6 | microJy            |5.23E+13|  8.22E-05|+/-2.76E-05|Jy|2007ApJS..171..353S|uncertainty|   5.731   microns   | Broad-band measurement|03 52 51.6 -27 49 22.61 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
4|8.0 microns (IRAC)  | 79.3      |+/-26.5 | microJy            |3.81E+13|  7.93E-05|+/-2.65E-05|Jy|2007ApJS..171..353S|uncertainty|   7.872   microns   | Broad-band measurement|03 52 51.6 -27 49 22.61 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
5|24 microns (MIPS)   | 321.0     |+/-60.7 | microJy            |1.27E+13|  3.21E-04|+/-6.07E-05|Jy|2007ApJS..171..353S|uncertainty|   23.68   microns   | Broad-band measurement|03 52 51.6 -27 49 22.61 (J2000)| Flux in fixed aperture|13" diameter aperture                   |From reprocessed raw data
6|70 microns (MIPS)   ||<1040      | microJy            |4.20E+12||1.04E-03|Jy|2007ApJS..171..353S|3 sigma|   71.42   microns   | Broad-band measurement|03 52 51.6 -27 49 22.61 (J2000)| Flux in fixed aperture|35" diameter aperture                   |From reprocessed raw data
7|160 microns (MIPS)  ||<88800     | microJy            |1.92E+12||8.88E-02|Jy|2007ApJS..171..353S|3 sigma|   155.9   microns   | Broad-band measurement|03 52 51.6 -27 49 22.61 (J2000)| Flux in fixed aperture|50" diameter aperture                   |From reprocessed raw data
8|4.85 GHz            | 86        |+/-11   |milliJy             |4.85E+09|  8.60E-02|+/-1.10E-02|Jy|1994ApJS...90..179G|rms noise|4.85       GHz       | Broad-band measurement|035249.2 -274948 (J2000)| Modelled datum|                                        |From new raw data; Corrected for contaminating sources
9|1.4GHz              | 350.3     |+/-10.5 |milliJy             |1.40E+09|  3.50E-01|+/-1.05E-02|Jy|1998AJ....115.1693C|uncertainty|    1.40   GHz       | Broad-band measurement|03 52 51.63 -27 49 23.0 (J2000)| Flux integrated from map|                                        |From new raw data
10|408 MHz             | 1.24      |+/-0.08 |Jy                  |4.08E+08|  1.24E+00|+/-8.00E-02|Jy|1981MNRAS.194..693L|rms noise|408        MHz       | Broad-band measurement|035048.1 -275812 (B1950)| Modelled datum|                                        |From new raw data; Corrected for contaminating sources
11|365 MHz (Texas)     | 1.636     |+/-0.069|Jy                  |3.65E+08|  1.64E+00|+/-6.90E-02|Jy|1996AJ....111.1945D|internal error|365        MHz       | Broad-band measurement; obtained by interpolation over frequency|035047.885 -275814.51 (B1950)| Integrated from scans|Model:D;MFlag:+;EFlag:+;LFlag:+.        |From new raw data
12|74 MHz (VLA)        | 4.15      |+/-0.43 | Jy                 |7.38E+07|  4.15E+00|+/-4.30E-01|Jy|2007AJ....134.1245C|rms uncertainty|    73.8   MHz       | Broad-band measurement|03 52 51.47 -27 49 24.3 (J2000)| Flux integrated from map|Corrected for clean bias                |From new raw data
