
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-02-19T12:27:01PST



Photometric Data for H-ATLASJ142413.9+023040

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|250 microns Herschel| 115       |+/-19   |milliJy             |1.20E+12|  1.15-01|+/-1.9E-02|Jy|2010A&A...518L..35I|uncertainty|       250 microns   | Broad-band measurement| | Flux integrated from map|                                        |From new raw data
2|350 microns Herschel| 192       |+/-30   |milliJy             |8.57E+11|  1.92E-01|+/-3.0E-02|Jy|2010A&A...518L..35I|uncertainty|       350 microns   | Broad-band measurement| | Flux integrated from map|                                        |From new raw data
3|500 microns Herschel| 204       |+/-32   |milliJy             |6.00E+11|  2.04-01|+/-3.2E-02|Jy|2010A&A...518L..35I|uncertainty|       500 microns   | Broad-band measurement| | Flux integrated from map|                                        |From new raw data
4|870 microns (APEX)  | 102       |+/-8.8  |milliJy             |3.45E+11|  1.02E-01|+/-8.8E-03|Jy|2010Natur.464..733S|uncertainty|       870 microns   | Broad-band measurement|21 35 11.6 -01 02 52.0 (J2000)| Flux in fixed aperture|                                        |From new raw data
5|880 microns (SMA)   | 90       |+/-5   |milliJy               |3.41E+11|  0.9E-01|+/-0.05E-02|Jy|2010Natur.464..733S|uncertainty|       434 microns   | Broad-band measurement|21 35 11.6 -01 02 52.0 (J2000)| Flux in fixed aperture|                                        |From new raw data
6|1.2 mm (MAMBO)      | 36        |+/-2    |milliJy             |2.50E+11|  3.60E-02|+/-2.00E-03|Jy|2010A&A...522L...4L|uncertainty|       1.2 mm        | Broad-band measurement|18 42 22.5 +59 38 30 (J2000)| Flux integrated from map|                                        |From new raw data
7|2.0 mm (PdBI)      | 9.7       |+/-0.9  |milliJy             |1.54E+11|  9.7E-03|+/-0.9E-04|Jy|2010Natur.464..733S|uncertainty|       2.8 microns   | Broad-band measurement|21 35 11.6 -01 02 52.0 (J2000)| Flux in fixed aperture|                                        |From new raw data
8|2.8 mm (PdBI)      | 1.8       |+/-0.3  |milliJy             |1.07E+11|  1.80E-03|+/-3.00E-04|Jy|2010Natur.464..733S|uncertainty|       2.8 microns   | Broad-band measurement|21 35 11.6 -01 02 52.0 (J2000)| Flux in fixed aperture|                                        |From new raw data
9|3.0mm (PdBI)       | 1.6       |+/-0.2  |milliJy             |9.99E+10|1.6E-03 |+/-0.2E-03|Jy|1995ApJ...450..559B|rms noise|1.4        GHz       | Broad-band measurement; synthetic band|120046.812 +300414.82 (J2000)| Peak flux|                                        |From new raw data; Corrected for contaminating sources
10|3.3mm (PdBI)       | 1.2       |+/-0.1   |milliJy             |9.11E+10|1.2E-03 |+/-0.1E-03|Jy|1995ApJ...450..559B|rms noise|1.4        GHz       | Broad-band measurement; synthetic band|120046.812 +300414.82 (J2000)| Peak flux|                                        |From new raw data; Corrected for contaminating sources
