
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-06-10T01:56:41PDT



Photometric Data for GOODS J123653.37+621140.0

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|4.0-8 keV (Chandra) ||<0.19E-15  |ergs cm^-2^ s^-1^   |1.45E+18||1.31E-11|Jy|2003AJ....126..539A|3 sigma|       6   keV       | Broad-band measurement|12 36 53.37 +62 11 39.6 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
2|4-8 keV (Chandra)   ||<0.17E-15  |erg cm^-2^ s^-1^    |1.45E+18||1.17E-11|Jy|2001AJ....122.2810B|3rms uncertainty reported|       6   keV       | Broad-band measurement|12 36 53.41 +62 11 39.6 (J2000)| Flux in fixed aperture|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
3|2-8 keV (Chandra)   ||<0.15E-15  |erg cm^-2^ s^-1^    |1.21E+18||1.24E-11|Jy|2001AJ....122.2810B|3rms uncertainty reported|       5   keV       | Broad-band measurement|12 36 53.41 +62 11 39.6 (J2000)| Flux in fixed aperture|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
4|2.0-8 keV (Chandra) ||<0.13E-15  |ergs cm^-2^ s^-1^   |1.21E+18||1.08E-11|Jy|2003AJ....126..539A|3 sigma|       5   keV       | Broad-band measurement|12 36 53.37 +62 11 39.6 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
5|0.5-8 keV (Chandra) | 0.22E-15  |+/-4   %|erg cm^-2^ s^-1^    |1.03E+18|  2.14E-11|+/-8.54E-13|Jy|2001AJ....122.2810B|estimated error|    4.25   keV       | Broad-band measurement|12 36 53.41 +62 11 39.6 (J2000)| Flux in fixed aperture|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
6|0.5-8 keV (Chandra) | 0.21E-15  ||ergs cm^-2^ s^-1^   |1.03E+18|  2.04E-11||Jy|2003AJ....126..539A|no uncertainty reported|    4.25   keV       | Broad-band measurement|12 36 53.37 +62 11 39.6 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
7|2.0-4 keV (Chandra) ||<0.11E-15  |ergs cm^-2^ s^-1^   |7.25E+17||1.52E-11|Jy|2003AJ....126..539A|3 sigma|       3   keV       | Broad-band measurement|12 36 53.37 +62 11 39.6 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
8|1.0-2 keV (Chandra) | 0.07E-15  ||ergs cm^-2^ s^-1^   |3.63E+17|  1.93E-11||Jy|2003AJ....126..539A|no uncertainty reported|     1.5   keV       | Broad-band measurement|12 36 53.37 +62 11 39.6 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
9|0.5-2 keV (Chandra) | 0.11E-15  ||ergs cm^-2^ s^-1^   |3.02E+17|  3.64E-11||Jy|2003AJ....126..539A|no uncertainty reported|    1.25   keV       | Broad-band measurement|12 36 53.37 +62 11 39.6 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
10|0.5-2 keV (Chandra) | 0.09E-15  |+/-4   %|erg cm^-2^ s^-1^    |3.02E+17|  2.98E-11|+/-1.19E-12|Jy|2001AJ....122.2810B|estimated error|    1.25   keV       | Broad-band measurement|12 36 53.41 +62 11 39.6 (J2000)| Flux in fixed aperture|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
11|0.5-1 keV (Chandra) | 0.05E-15  ||ergs cm^-2^ s^-1^   |1.81E+17|  2.76E-11||Jy|2003AJ....126..539A|no uncertainty reported|    0.75   keV       | Broad-band measurement|12 36 53.37 +62 11 39.6 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
12|U (KPNO) AB         | 22.78     ||mag                 |8.44E+14|  2.81E-06||Jy|2006ApJ...653.1004R|no uncertainty reported|    3550   A         | Broad-band measurement|123653.46 +621140.0 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data; derived from aflux in a different band and a color
13|U (KPNO) AB         | 23.4      || mag                |8.22E+14|  1.59E-06||Jy|2004AJ....127.3137C|no uncertainty reported| 3647.65   A         | Broad-band measurement|189.222382 +62.19444 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
14|B (HST/ACS) AB      | 23.298    ||mag                 |6.98E+14|  1.74E-06||Jy|2007ApJ...660...81M|no uncertainty reported|    4297   A         | Broad-band measurement|12 36 53.383 +62 11 39.57 (J2000)| Flux integrated from map|                                        |From reprocessed raw data; Corrected for contaminatingsources
15|B (SUBARU) AB       | 23.32     ||mag                 |6.77E+14|  1.71E-06||Jy|2006ApJ...653.1027W|no uncertainty reported| 4427.60   A         | Broad-band measurement|189.222429 62.194325 (J2000)| Flux in fixed aperture|3" diameter aperture                    |Averaged from previously published data
16|B (Subaru) AB       | 23.3      || mag                |6.77E+14|  1.74E-06||Jy|2004AJ....127.3137C|no uncertainty reported| 4427.60   A         | Broad-band measurement|189.222382 +62.19444 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
17|G (KECK) AB         | 22.59     ||mag                 |6.27E+14|  3.34E-06||Jy|2006ApJ...653.1004R|no uncertainty reported|    4780   A         | Broad-band measurement|123653.46 +621140.0 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data; derived from aflux in a different band and a color
18|V (Subaru) AB       | 23.2      || mag                |5.48E+14|  1.91E-06||Jy|2004AJ....127.3137C|no uncertainty reported| 5471.22   A         | Broad-band measurement|189.222382 +62.19444 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
19|V (HST/ACS) AB      | 22.915    ||mag                 |5.08E+14|  2.48E-06||Jy|2007ApJ...660...81M|no uncertainty reported|    5907   A         | Broad-band measurement|12 36 53.383 +62 11 39.57 (J2000)| Flux integrated from map|                                        |From reprocessed raw data; Corrected for contaminatingsources
20|R (Keck II) AB      | 23.05     || mag                |4.62E+14|  2.19E-06||Jy|2004AJ....127.3121W|no uncertainty reported|   648.7   A         | Broad-band measurement|12 36 53.383 +62 11 39.57 (J2000)| Total flux|                                        |From new raw data
21|R (SUBARU) AB       | 22.93     ||mag                 |4.59E+14|  2.44E-06||Jy|2006ApJ...653.1027W|no uncertainty reported| 6534.16   A         | Broad-band measurement|189.222429 62.194325 (J2000)| Flux in fixed aperture|3" diameter aperture                    |Averaged from previously published data
22|R (Subaru) AB       | 22.9      || mag                |4.59E+14|  2.51E-06||Jy|2004AJ....127.3137C|no uncertainty reported| 6534.16   A         | Broad-band measurement|189.222382 +62.19444 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
23|R (SUBARU) AB       | 22.93     ||mag                 |4.58E+14|  2.44E-06||Jy|2007MNRAS.377..203G|no uncertainty reported|    6550   A         | Broad-band measurement|12 36 53.37 +62 11 39.6 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
24|R (KECK) AB         | 22.31     ||mag                 |4.39E+14|  4.33E-06||Jy|2006ApJ...653.1004R|no uncertainty reported|    6830   A         | Broad-band measurement|123653.46 +621140.0 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data
25|i (HST/ACS) AB      | 22.410    ||mag                 |3.86E+14|  3.95E-06||Jy|2007ApJ...660...81M|no uncertainty reported|    7764   A         | Broad-band measurement|12 36 53.383 +62 11 39.57 (J2000)| Flux integrated from map|                                        |From reprocessed raw data; Corrected for contaminatingsources
26|I (SUBARU) AB       | 22.51     ||mag                 |3.76E+14|  3.60E-06||Jy|2006ApJ...653.1027W|no uncertainty reported| 7975.89   A         | Broad-band measurement|189.222429 62.194325 (J2000)| Flux in fixed aperture|3" diameter aperture                    |Averaged from previously published data
27|I (Subaru) AB       | 22.5      || mag                |3.76E+14|  3.63E-06||Jy|2004AJ....127.3137C|no uncertainty reported| 7975.89   A         | Broad-band measurement|189.222382 +62.19444 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
28|z' (Subaru) AB      | 22.1      || mag                |3.31E+14|  5.25E-06||Jy|2004AJ....127.3137C|no uncertainty reported| 9069.21   A         | Broad-band measurement|189.222382 +62.19444 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
29|z (HST/ACS) AB      | 21.954    ||mag                 |3.17E+14|  6.00E-06||Jy|2007ApJ...660...81M|no uncertainty reported|    9445   A         | Broad-band measurement|12 36 53.383 +62 11 39.57 (J2000)| Flux integrated from map|                                        |From reprocessed raw data; Corrected for contaminatingsources
30|J (WIRC) AB         | 21.46     ||mag                 |2.40E+14|  9.46E-06||Jy|2006ApJ...653.1004R|no uncertainty reported|   1.250   microns   | Broad-band measurement|123653.46 +621140.0 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data
31|HK' (QUIRC) AB      | 21.11     |+/-0.06 |mag                 |1.58E+14|  1.31E-05|+/-7.22E-07|Jy|2006ApJ...653.1027W|uncertainty|18947.38   A         | Broad-band measurement|189.222429 62.194325 (J2000)| Flux in fixed aperture|3" diameter aperture                    |Averaged from previously published data
32|HK' (UH) AB         | 21.1      || mag                |1.58E+14|  1.32E-05||Jy|2004AJ....127.3137C|no uncertainty reported|18947.38   A         | Broad-band measurement|189.222382 +62.19444 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
33|K_s (Hale/WIRC) AB  | 20.47     ||mag                 |1.39E+14|  2.36E-05||Jy|2005ApJ...633..748R|no uncertainty reported|   2.150   microns   | Broad-band measurement|12 36 53.46 +62 11 40.0 (J2000)| Flux in fixed aperture|                                        |From new raw data
34|K_s (WIRC) AB       | 20.47     ||mag                 |1.39E+14|  2.36E-05||Jy|2006ApJ...653.1004R|no uncertainty reported|   2.150   microns   | Broad-band measurement|123653.46 +621140.0 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data
35|3.6 microns IRAC AB | 20.38     |+/-0.07 |mag                 |8.44E+13|  2.56E-05|+/-1.65E-06|Jy|2006ApJ...653.1004R|uncertainty|   3.550   microns   | Broad-band measurement|123653.46 +621140.0 (J2000)| Flux integrated from map|                                        |From new raw data
36|3.6 microns (IRAC)  | 33.50     |+/-0.06 |microJy             |8.44E+13|  3.35E-05|+/-6.00E-08|Jy|2007MNRAS.377..203G|uncertainty|   3.550   microns   | Broad-band measurement|12 36 53.37 +62 11 39.6 (J2000)| Corrected to total flux from single aperture measurement|                                        |From reprocessed raw data
37|3.6 microns (IRAC)  | 33.60     |+/-1.68 |microJy             |8.44E+13|  3.36E-05|+/-1.68E-06|Jy|2011AJ....141....1T|rms uncertainty|     3.550 microns   | Broad-band measurement|189.222397 62.194351 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
38|4.5 microns (IRAC)  | 36.86     |+/-0.09 |microJy             |6.67E+13|  3.69E-05|+/-9.00E-08|Jy|2007MNRAS.377..203G|uncertainty|   4.493   microns   | Broad-band measurement|12 36 53.37 +62 11 39.6 (J2000)| Corrected to total flux from single aperture measurement|                                        |From reprocessed raw data
39|4.5 microns IRAC AB | 20.29     |+/-0.07 |mag                 |6.67E+13|  2.78E-05|+/-1.79E-06|Jy|2006ApJ...653.1004R|uncertainty|   4.493   microns   | Broad-band measurement|123653.46 +621140.0 (J2000)| Flux integrated from map|                                        |From new raw data
40|4.5 microns (IRAC)  | 36.40     |+/-1.82 |microJy             |6.67E+13|  3.64E-05|+/-1.82E-06|Jy|2011AJ....141....1T|rms uncertainty|     4.493 microns   | Broad-band measurement|189.222397 62.194351 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
41|5.8 microns IRAC AB | 20.48     |+/-0.07 |mag                 |5.23E+13|  2.33E-05|+/-1.50E-06|Jy|2006ApJ...653.1004R|uncertainty|   5.731   microns   | Broad-band measurement|123653.46 +621140.0 (J2000)| Flux integrated from map|                                        |From new raw data
42|5.8 microns (IRAC)  | 30.47     |+/-0.48 |microJy             |5.23E+13|  3.05E-05|+/-4.80E-07|Jy|2007MNRAS.377..203G|uncertainty|   5.731   microns   | Broad-band measurement|12 36 53.37 +62 11 39.6 (J2000)| Corrected to total flux from single aperture measurement|                                        |From reprocessed raw data
43|5.8 microns (IRAC)  | 28.90     |+/-1.49 |microJy             |5.23E+13|  2.89E-05|+/-1.49E-06|Jy|2011AJ....141....1T|rms uncertainty|     5.731 microns   | Broad-band measurement|189.222397 62.194351 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
44|8.0 microns IRAC AB | 20.02     |+/-0.07 |mag                 |3.81E+13|  3.56E-05|+/-2.30E-06|Jy|2006ApJ...653.1004R|uncertainty|   7.872   microns   | Broad-band measurement|123653.46 +621140.0 (J2000)| Flux integrated from map|                                        |From new raw data
45|8.0 microns (IRAC)  | 42.51     |+/-0.50 |microJy             |3.81E+13|  4.25E-05|+/-5.00E-07|Jy|2007MNRAS.377..203G|uncertainty|   7.872   microns   | Broad-band measurement|12 36 53.37 +62 11 39.6 (J2000)| Corrected to total flux from single aperture measurement|                                        |From reprocessed raw data
46|8.0 microns (IRAC)  | 41.80     |+/-2.13 |microJy             |3.81E+13|  4.18E-05|+/-2.13E-06|Jy|2011AJ....141....1T|rms uncertainty|     7.872 microns   | Broad-band measurement|189.222397 62.194351 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
47|11 microns (AKARI)  | 57.0      |+/-15   | microJy            |2.73E+13|  5.70E-05|+/-1.50E-05|Jy|2009MNRAS.394..375N|uncertainty|        11 microns   | Broad-band measurement|12 36 53.37 +62 11 39.97 (J2000)| Flux integrated from map|                                        |From new raw data
48|ISOCAM 15 microns   | 0.1382    |+/-0.1  |milliJy             |2.07E+13|  1.38E-04|+/-1.00E-04|Jy|1997MNRAS.289..465G|estimated error|14.5       microns   | Broad-band measurement|123653.05 +621116.9 (J2000)| Flux integrated from map|                                        |From new raw data
49|15 microns (ISOCAM) | 180       |+/-36   |microJy             |2.00E+13|  1.80E-04|+/-3.60E-05|Jy|2006A&A...451...57M|68% confidence|    15.0   microns   | Broad-band measurement|189.2223816 62.1944351 (J2000)| Flux integrated from map|                                        |Averaged from previously published data
50|16 microns (IRS)    | 436.6     |+/-10.0 |microJy             |1.90E+13|  4.37E-04|+/-1.00E-05|Jy|2011AJ....141....1T|rms uncertainty|      15.8 microns   | Broad-band measurement|189.222397 62.194351 (J2000)| From fitting to map|                                        |From new raw data
51|18 microns (AKARI)  | 393       |+/-33   | microJy            |1.67E+13|  3.93E-04|+/-3.30E-05|Jy|2009MNRAS.394..375N|uncertainty|        18 microns   | Broad-band measurement|12 36 53.37 +62 11 39.97 (J2000)| Flux integrated from map|                                        |From new raw data
52|24 microns (MIPS)   | 322       |+/-6    |microJy             |1.27E+13|  3.22E-04|+/-6.00E-06|Jy|2006A&A...451...57M|68% confidence|   23.68   microns   | Broad-band measurement|189.2223816 62.1944351 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
53|24 microns (MIPS)   | 303.2     |+/-17.6 |microJy             |1.27E+13|  3.03E-04|+/-1.76E-05|Jy|2006ApJ...653.1004R|uncertainty|   23.68   microns   | Broad-band measurement|123653.46 +621140.0 (J2000)| Flux integrated from map|                                        |From new raw data
54|24 microns (MIPS)   | 319.76    |+/-4.90 |microJy             |1.27E+13|  3.20E-04|+/-4.90E-06|Jy|2007MNRAS.377..203G|uncertainty|   23.68   microns   | Broad-band measurement|12 36 53.37 +62 11 39.6 (J2000)| Corrected to total flux from single aperture measurement|                                        |From reprocessed raw data
55|24 microns (MIPS)   | 336.0     |+/-7.5  |microJy             |1.27E+13|  3.36E-04|+/-7.50E-06|Jy|2011AJ....141....1T|rms uncertainty|     23.68 microns   | Broad-band measurement|189.222397 62.194351 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
56|24 microns (Spitzer)| 322       |+/-6    |microJy             |1.27E+13|  3.22E-04|+/-6.00E-06|Jy|2011ApJ...726...93R|uncertainty|     23.68 microns   | Broad-band measurement|12 36 53.37 +62 11 39.6 (J2000)| Not reported in paper|                                        |Averaged from previously published data
60|24 microns (MIPS)   | 339.2     |+/-4.5  |microJy             |1.27E+13|  3.39E-04|+/-4.50E-06|Jy|2011A&A...528A..35M|uncertainty|     23.68 microns   | Broad-band measurement|12 36 53.38 +62 11 39.60 (J2000)| Flux integrated from map|                                        |From new raw data
57|70 microns (Spitzer)| 6.6       |+/-0.4  | milliJy            |4.20E+12|  6.60E-03|+/-4.00E-04|Jy|2009MNRAS.399..121C|uncertainty|     71.42 microns   | Broad-band measurement|123653.37 +621139.6 (J2000)| Flux integrated from map|                                        |From reprocessed raw data
62|70 microns (MIPS)   | 7.6       |+/-0.3  |milliJy             |4.20E+12|  7.60E-03|+/-3.00E-04|Jy|2011A&A...528A..35M|uncertainty|     71.42 microns   | Broad-band measurement|12 36 53.38 +62 11 39.60 (J2000)| Flux integrated from map|                                        |From new raw data
58|850 microns (SCUBA) ||<1.4       | milliJy            |3.53E+11||1.40E-03|Jy|2009MNRAS.399..121C|2 sigma|       850 microns   | Broad-band measurement|123653.37 +621139.6 (J2000)| Flux integrated from map|                                        |From new raw data
58|850 microns (SCUBA) ||<1.8       | milliJy            |3.53E+11||1.80E-03|Jy|2009MNRAS.399..121C|3 sigma|       850 microns   | Broad-band measurement|123653.37 +621139.6 (J2000)| Flux integrated from map|                                        |From new raw data
4|1200 microns (MAMBO)|           |<1.1    |mJy             |2.50E+11|        |1.1E-03|Jy|2004MNRAS.354..779G|3rms uncertainty|      1200 microns   | Broad-band measurement|16 36 55.9 +40 59 12 (J2000)| Flux integrated from map|S/N = 3.66                              |From new raw data
59|8.5 GHz             | 12.60     ||microJy             |8.50E+09|  1.26E-05||Jy|1998AJ....116.1039R|no uncertainty reported|8.5        GHz       | Broad-band measurement; peak value reported; synthetic band|123653.348 +621139.54 (J2000)| Flux integrated from map; Pointing and beam filling|                                        |From new raw data; Corrected for contaminating sources
60|8.5 GHz             | 12.60     ||microJy             |8.50E+09|  1.26E-05||Jy|1998AJ....116.1039R|no uncertainty reported|8.5        GHz       | Broad-band measurement; broad-band flux derived by integration over spectrum; synthetic band|123653.348 +621139.54 (J2000)| Flux integrated from map; Pointing and beam filling|                                        |From new raw data; Corrected for contaminating sources
61|8.4 GHz             | 15        |+/-3    |uJy                 |8.40E+09|  1.50E-05|+/-3.00E-06|Jy|1997ApJ...475L...5F|estimated error| 8.4       GHz       | Broad-band measurement|123653.35 +621139.7 (J2000)| Flux integrated from map; Beam filling or dilution corrected|                                        |From new raw data
62|1.4 GHz (VLA)       | 62        |+/-6    | microJy            |1.40E+09|  6.20E-05|+/-6.00E-06|Jy|2006MNRAS.371..963B|1 sigma|       1.4 GHz       | Broad-band measurement|12 36 53.374 +62 11 39.68 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
63|1.4 GHz (VLA)       | 73.97     ||microJy             |1.40E+09|  7.40E-05||Jy|2006A&A...451...57M|no uncertainty reported|     1.4   GHz       | Broad-band measurement|189.2223816 62.1944351 (J2000)| Flux integrated from map|                                        |From new raw data
64|1.4 GHz (VLA)       | 66        ||microJy             |1.40E+09|  6.60E-05||Jy|2005MNRAS.358.1159M|no uncertainty reported|     1.4   GHz       | Broad-band measurement|12 36 53.3629 +62 11 39.647 (J2000)| Flux integrated from map|                                        |From new raw data
65|1.4 GHz (MERLIN)    | 86.7      |+/-8.3  | microJy            |1.40E+09|  8.67E-05|+/-8.30E-06|Jy|2009MNRAS.399..121C|uncertainty|       1.4 GHz       | Broad-band measurement|123653.37 +621139.6 (J2000)| Flux integrated from map|                                        |From new raw data
66|1.4 GHz             | 65.7      |+/-8.2  |microJy             |1.40E+09|  6.57E-05|+/-8.20E-06|Jy|2000ApJ...533..611R|1 sigma|1.4        GHz       | Broad-band measurement; broad-band flux derived by integration over spectrum; synthetic band|123653.402 +621139.61 (J2000)| Flux integrated from map; Pointing and beam filling|                                        |From new raw data; Corrected for contaminating sources
67|1.4 GHz (VLA)       | 84.2      |+/-8.9  |microJy             |1.40E+09|  8.42E-05|+/-8.90E-06|Jy|2010ApJS..188..178M|uncertainty|       1.4 GHz       | Broad-band measurement|12 36 53.35 +62 11 39.7 (J2000)| Total flux; Beam filling or dilution corrected|Major=1.0"; Minor=0.5"; PA=32 deg       |From new raw data
