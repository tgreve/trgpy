
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-06-16T17:17:01PDT



Photometric Data for [HB89] 2343+125:BX0610

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|G (WHT)             | 23.92     ||mag                 |6.38E+14|  9.82E-07||Jy|2006ApJ...647..128E|no uncertainty reported|    0.47   microns   | Broad-band measurement|| Flux in fixed aperture|                                        |Averaged from previously published data
2|H{beta} (VLT)       | 0.61E-16  |+/-0.08E-16|erg/s/cm^2^         |6.17E+14|  6.10E+06|+/-8.00E+05|Jy-Hz|2009ApJ...699.1660L|uncertainty|      4861 A         | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|                                        |From new raw data
3|H{alpha} (Keck II)  | 8.1E-17   |+/-0.4E-17|erg s^-1^ cm^-2^    |4.57E+14|  8.10E+06|+/-4.00E+05|Jy-Hz|2006ApJ...646..107E|uncertainty|    6563   A         | Line measurement; flux integrated over line; lines measured in emission|23 46 09.43 +12 49 19.21 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
4|H{alpha} (VLT)      | 30.5E-17  |+/-1.3E-17|erg/s/cm^2^         |4.57E+14|  3.05E+07|+/-1.30E+06|Jy-Hz|2009ApJ...706.1364F|uncertainty|      6563 A         | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|                                        |From new raw data
5|[S II] 6716 (VLT)   | 1.7E-16   |+/-0.1E-16|erg/s/cm^2^         |4.46E+14|  1.70E+07|+/-1.00E+06|Jy-Hz|2009ApJ...699.1660L|uncertainty|      6716 A         | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|                                        |From new raw data
6|[S II] 6731 (VLT)   | 1.5E-16   |+/-0.1E-16|erg/s/cm^2^         |4.45E+14|  1.50E+07|+/-1.00E+06|Jy-Hz|2009ApJ...699.1660L|uncertainty|      6731 A         | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|                                        |From new raw data
7|J (Hale/WIRC)       | 21.45     ||mag                 |2.40E+14|  4.10E-06||Jy|2006ApJ...646..107E|no uncertainty reported|    1.25   microns   | Broad-band measurement|23 46 09.43 +12 49 19.21 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data; derived from aflux in a different band and a color
8|F160W (HST) AB      | 22.09     |+/-0.06 |mag                 |1.87E+14|  5.30E-06|+/-2.93E-07|Jy|2011ApJ...731...65F|uncertainty|     1.603 microns   | Broad-band measurement|| Flux in fixed aperture|                                        |From new raw data
9|K_s (Hale/WIRC)     | 19.21     ||mag                 |1.39E+14|  1.39E-05||Jy|2006ApJ...646..107E|no uncertainty reported|    2.15   microns   | Broad-band measurement|23 46 09.43 +12 49 19.21 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data
10|CO(3-2) (PdBI)      ||<0.08      |Jy km/s             |3.46E+11|  3.42E+05|2.88E+04|Jy-Hz|2010Natur.463..781T|3 sigma|   345.998 GHz       | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|                                        |From new raw data
