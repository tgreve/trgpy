
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-06-16T17:07:52PDT



Photometric Data for CXOU J170054.48+641623.8

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|U_n (WHT) AB        | 26.38     |+/-0.33 |mag                 |8.33E+14|  1.02E-07|+/-3.06E-08|Jy|2005ApJ...626..698S|estimated error|    0.36   microns   | Broad-band measurement|17 00 54.542 64 16 24.760 (J2000)| Flux integrated from map|                                        |From new raw data; derived from a flux in a different bandand a color
2|G (WHT) AB          | 24.88     |+/-0.18 |mag                 |6.38E+14|  4.05E-07|+/-6.86E-08|Jy|2005ApJ...626..698S|estimated error|    0.47   microns   | Broad-band measurement|17 00 54.542 64 16 24.760 (J2000)| Flux integrated from map|                                        |From new raw data; derived from a flux in a different bandand a color
3|G (WHT)             | 24.88     ||mag                 |6.38E+14|  4.05E-07||Jy|2006ApJ...647..128E|no uncertainty reported|    0.47   microns   | Broad-band measurement|| Flux in fixed aperture|                                        |Averaged from previously published data
4|H{alpha} (Keck II)  | 12.9E-17  |+/-1.4E-17|erg s^-1^ cm^-2^    |4.57E+14|  1.29E+07|+/-1.40E+06|Jy-Hz|2006ApJ...646..107E|uncertainty|    6563   A         | Line measurement; flux integrated over line; lines measured in emission|17 00 54.54 +64 16 24.76 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
5|R (WHT) AB          | 24.56     |+/-0.16 |mag                 |4.41E+14|  5.44E-07|+/-8.02E-08|Jy|2005ApJ...626..698S|estimated error|    0.68   microns   | Broad-band measurement|17 00 54.542 64 16 24.760 (J2000)| Flux integrated from map|                                        |From new raw data
6|J (Hale/WIRC)       | 19.90     ||mag                 |2.40E+14|  1.71E-05||Jy|2006ApJ...646..107E|no uncertainty reported|    1.25   microns   | Broad-band measurement|17 00 54.54 +64 16 24.76 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data; derived from aflux in a different band and a color
7|K_s (Hale/WIRC)     | 19.90     ||mag                 |1.39E+14|  7.35E-06||Jy|2006ApJ...646..107E|no uncertainty reported|    2.15   microns   | Broad-band measurement|17 00 54.54 +64 16 24.76 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data
8|K_s (P200) AB       | 21.64     |+/-0.19 |mag                 |1.39E+14|  8.02E-06|+/-1.43E-06|Jy|2005ApJ...626..698S|estimated error|    2.15   microns   | Broad-band measurement|17 00 54.542 64 16 24.760 (J2000)| Flux integrated from map|                                        |From new raw data; derived from a flux in a different bandand a color
9|4.5 microns IRAC AB | 20.51     |+/-0.10 |mag                 |6.66E+13|  2.27E-05|+/-2.09E-06|Jy|2005ApJ...626..698S|estimated error|     4.5   microns   | Broad-band measurement|17 00 54.542 64 16 24.760 (J2000)| Flux integrated from map|                                        |From new raw data
10|8.0 microns IRAC AB | 18.51     |+/-0.10 |mag                 |3.75E+13|  1.43E-04|+/-1.32E-05|Jy|2005ApJ...626..698S|estimated error|     8.0   microns   | Broad-band measurement|17 00 54.542 64 16 24.760 (J2000)| Flux integrated from map|                                        |From new raw data
11|CO(3-2) (PdBI)      ||<0.08      |Jy km/s             |3.46E+11|  2.07E+05|2.76E+04|Jy-Hz|2010Natur.463..781T|3 sigma|   345.998 GHz       | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|                                        |From new raw data
