
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-04-04T08:30:18PDT



Photometric Data for SMM J163541.2+661144

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|450 microns (SCUBA) | |<59.4      |milliJy             |6.66E+11| |5.94E-02|Jy|2006MNRAS.368..487K|3rms uncertainty reported|     450   microns   | Broad-band measurement|163541.2 +661144 (J2000)| Flux integrated from map|                                        |From new raw data
2|450 microns (SCUBA) | 53.4      |+/-16.0 | milliJy            |6.66E+11|  5.34E-02|+/-1.60E-02|Jy|2008MNRAS.384.1611K|rms uncertainty|       450 microns   | Broad-band measurement|163541.2 +661144 (J2000)| Flux integrated from map|S/N = 3.5                               |From new raw data
3|850 microns (SCUBA) | 10.4      |+/-1.4  | milliJy            |3.53E+11|  1.04E-02|+/-1.40E-03|Jy|2008MNRAS.384.1611K|rms uncertainty|       850 microns   | Broad-band measurement|163541.2 +661144 (J2000)| Flux integrated from map|S/N = 7.5                               |From new raw data
4|850 microns (SCUBA) | 10.4      |+/-1.4  |milliJy             |3.53E+11|  1.04E-02|+/-1.40E-03|Jy|2006MNRAS.368..487K|uncertainty|     850   microns   | Broad-band measurement|163541.2 +661144 (J2000)| Flux integrated from map|                                        |From new raw data
5|CO(3-2) (IRAM)      | 1.0       |+/-0.1  | Jy km/s            |3.46E+11|  1.91E-07|+/-1.91E-08|Jy|2009A&A...496...45K|uncertainty|   345.796 GHz       | Line measurement; flux integrated over line; lines measured in emission|16 35 40.86 +66 11 44.4 (J2000)| Flux integrated from map|                                        |From new raw data
6|CO(3-2) (IRAM)      | 0.3       |+/-0.1  | Jy km/s            |3.46E+11|  5.70E-08|+/-1.90E-08|Jy|2009A&A...496...45K|uncertainty|   345.796 GHz       | Line measurement; flux integrated over line; lines measured in emission|16 35 41.33 +66 11 46.4 (J2000)| Flux integrated from map|                                        |From new raw data
7|3 mm (IRAM)         | |<0.6       | milliJy            |9.99E+10| |6.00E-04|Jy|2009A&A...496...45K|3rms uncertainty|         3 mm        | Broad-band measurement|16 35 41.33 +66 11 46.4 (J2000)| Flux integrated from map|                                        |From new raw data
