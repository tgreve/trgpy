
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-06-11T21:22:18PDT



Photometric Data for GOODS J123707.21+621408.1

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|4.0-8 keV (Chandra) | 0.60E-15  ||ergs cm^-2^ s^-1^   |1.45E+18|  4.14E-11||Jy|2003AJ....126..539A|no uncertainty reported|       6   keV       | Broad-band measurement|12 37 07.20 +62 14 07.9 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
2|4-8 keV (Chandra)   | 0.63E-15  |+/-4   %|erg cm^-2^ s^-1^    |1.45E+18|  4.34E-11|+/-1.74E-12|Jy|2001AJ....122.2810B|estimated error|       6   keV       | Broad-band measurement|12 37 07.23 +62 14 08.0 (J2000)| Flux in fixed aperture|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
3|2-10 keV (Chandra)  | 7.38E-16  ||erg/cm^2^/s         |1.45E+18|  5.09E-11||Jy|2010MNRAS.401.2763L|no uncertainty reported|      6.00 keV       | Broad-band measurement|189.279970 62.235370 (J2000)| Modelled datum|                                        |From reprocessed raw data; NED frequency assigned tomid-point of band in keV
4|2-8 keV (Chandra)   | 0.92E-15  |+/-4   %|erg cm^-2^ s^-1^    |1.21E+18|  7.60E-11|+/-3.04E-12|Jy|2001AJ....122.2810B|estimated error|       5   keV       | Broad-band measurement|12 37 07.23 +62 14 08.0 (J2000)| Flux in fixed aperture|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
5|2.0-8 keV (Chandra) | 0.91E-15  ||ergs cm^-2^ s^-1^   |1.21E+18|  7.53E-11||Jy|2003AJ....126..539A|no uncertainty reported|       5   keV       | Broad-band measurement|12 37 07.20 +62 14 07.9 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
6|0.5-8 keV (Chandra) | 1.00E-15  |+/-4   %|erg cm^-2^ s^-1^    |1.03E+18|  9.71E-11|+/-3.88E-12|Jy|2001AJ....122.2810B|estimated error|    4.25   keV       | Broad-band measurement|12 37 07.23 +62 14 08.0 (J2000)| Flux in fixed aperture|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
7|0.5-8 keV (Chandra) | 0.98E-15  ||ergs cm^-2^ s^-1^   |1.03E+18|  9.53E-11||Jy|2003AJ....126..539A|no uncertainty reported|    4.25   keV       | Broad-band measurement|12 37 07.20 +62 14 07.9 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
8|2.0-4 keV (Chandra) | 0.27E-15  ||ergs cm^-2^ s^-1^   |7.25E+17|  3.72E-11||Jy|2003AJ....126..539A|no uncertainty reported|       3   keV       | Broad-band measurement|12 37 07.20 +62 14 07.9 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
9|1.0-2 keV (Chandra) | 0.09E-15  ||ergs cm^-2^ s^-1^   |3.63E+17|  2.48E-11||Jy|2003AJ....126..539A|no uncertainty reported|     1.5   keV       | Broad-band measurement|12 37 07.20 +62 14 07.9 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
10|0.5-2 keV (Chandra) | 0.09E-15  ||ergs cm^-2^ s^-1^   |3.02E+17|  2.98E-11||Jy|2003AJ....126..539A|no uncertainty reported|    1.25   keV       | Broad-band measurement|12 37 07.20 +62 14 07.9 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
11|0.5-2 keV (Chandra) | 0.12E-15  |+/-4   %|erg cm^-2^ s^-1^    |3.02E+17|  3.97E-11|+/-1.59E-12|Jy|2001AJ....122.2810B|estimated error|    1.25   keV       | Broad-band measurement|12 37 07.23 +62 14 08.0 (J2000)| Flux in fixed aperture|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
12|0.5-1 keV (Chandra) ||<0.03E-15  |ergs cm^-2^ s^-1^   |1.81E+17||1.65E-11|Jy|2003AJ....126..539A|3 sigma|    0.75   keV       | Broad-band measurement|12 37 07.20 +62 14 07.9 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
13|U (KPNO/MOSAIC) AB  ||>27.8      |mag                 |8.44E+14||2.75E-08|Jy|2005ApJ...635..853B|2.5 sigma|    3552   A         | Broad-band measurement|123707.21 +621408.1 (J2000)| Flux in fixed aperture|3" aperture                             |Averaged new and previously published data
14|B (SUBARU) AB       | 26.77     |+/-0.27 |mag                 |6.81E+14|  7.11E-08|+/-1.77E-08|Jy|2005ApJ...635..853B|uncertainty|    4400   A         | Broad-band measurement|123707.21 +621408.1 (J2000)| Flux in fixed aperture|3" aperture                             |Averaged new and previously published data
15|V (SUBARU) AB       | 26.36     |+/-0.29 |mag                 |5.42E+14|  1.04E-07|+/-2.77E-08|Jy|2005ApJ...635..853B|uncertainty|    5530   A         | Broad-band measurement|123707.21 +621408.1 (J2000)| Flux in fixed aperture|3" aperture                             |Averaged new and previously published data
16|R (SUBARU) AB       | 25.63     |+/-0.14 |mag                 |4.68E+14|  2.03E-07|+/-2.62E-08|Jy|2005ApJ...635..853B|uncertainty|    6400   A         | Broad-band measurement|123707.21 +621408.1 (J2000)| Flux in fixed aperture|3" aperture                             |Averaged new and previously published data
17|H{alpha} (Keck)     | 1.6E-19   |+/-0.5E-19| W/m^2^             |4.57E+14|  1.60E+07|+/-5.00E+06|Jy-Hz|2004ApJ...617...64S|uncertainty|      6563 A         | Line measurement; flux integrated over line; lines measured in emission|123707.21 +621408.1 (J2000)| Flux integrated from map|                                        |From new raw data
18|I (SUBARU) AB       | 25.51     |+/-0.30 |mag                 |3.79E+14|  2.27E-07|+/-6.27E-08|Jy|2005ApJ...635..853B|uncertainty|    7900   A         | Broad-band measurement|123707.21 +621408.1 (J2000)| Flux in fixed aperture|3" aperture                             |Averaged new and previously published data
19|I (Cousins)         | 24.55     |+/-0.11 |mag                 |3.79E+14|  3.86E-07|+/-4.12E-08|Jy|2004ApJ...616...71S|1 sigma|    7900   A         | Broad-band measurement|| Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
20|z' (SUBARU) AB      | 24.69     |+/-0.19 |mag                 |3.30E+14|  4.83E-07|+/-8.45E-08|Jy|2005ApJ...635..853B|uncertainty|    9097   A         | Broad-band measurement|123707.21 +621408.1 (J2000)| Flux in fixed aperture|3" aperture                             |Averaged new and previously published data
21|J (Hale/WIRC) AB    ||>24.0      |mag                 |2.40E+14||9.12E-07|Jy|2005ApJ...635..853B|2.5 sigma|   1.250   microns   | Broad-band measurement|123707.21 +621408.1 (J2000)| Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
22|J (2MASS)           | 22.50     |+/-0.32 |mag                 |2.40E+14|  1.59E-06|+/-5.46E-07|Jy|2004ApJ...616...71S|1 sigma|    1.25   microns   | Broad-band measurement|| Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
23|K_s (Hale/WIRC) AB  | 21.87     ||mag                 |1.39E+14|  6.49E-06||Jy|2005ApJ...633..748R|no uncertainty reported|   2.150   microns   | Broad-band measurement|12 37 07.21 +62 14 08.1 (J2000)| Flux in fixed aperture|                                        |From new raw data
24|K_s_ (Hale/WIRC) AB | 21.86     |+/-0.11 |mag                 |1.39E+14|  6.55E-06|+/-6.63E-07|Jy|2005ApJ...635..853B|uncertainty|   2.150   microns   | Broad-band measurement|123707.21 +621408.1 (J2000)| Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
25|K_s_ (2MASS)        | 20.05     |+/-0.11 |mag                 |1.38E+14|  6.37E-06|+/-6.79E-07|Jy|2004ApJ...616...71S|1 sigma|    2.17   microns   | Broad-band measurement|| Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
26|3.6 microns IRAC AB | 20.68     |+/-0.10 |mag                 |8.44E+13|  1.94E-05|+/-1.79E-06|Jy|2005ApJ...635..853B|uncertainty|   3.550   microns   | Broad-band measurement|123707.21 +621408.1 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged new and previously published data
27|3.6 microns (IRAC)  | 18.7      |+/-2.2  |microJy             |8.44E+13|  1.87E-05|+/-2.20E-06|Jy|2009ApJ...699.1610H|uncertainty|     3.550 microns   | Broad-band measurement|12 37 07.20 +62 14 08.0 (J2000)| Flux in fixed aperture|                                        |From new raw data
28|4.5 microns IRAC AB | 20.33     |+/-0.08 |mag                 |6.67E+13|  2.68E-05|+/-1.97E-06|Jy|2005ApJ...635..853B|uncertainty|   4.493   microns   | Broad-band measurement|123707.21 +621408.1 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged new and previously published data
29|4.5 microns (IRAC)  | 24.2      |+/-2.5  |microJy             |6.67E+13|  2.42E-05|+/-2.50E-06|Jy|2009ApJ...699.1610H|uncertainty|     4.493 microns   | Broad-band measurement|12 37 07.20 +62 14 08.0 (J2000)| Flux in fixed aperture|                                        |From new raw data
30|5.8 microns IRAC AB | 20.02     |+/-0.14 |mag                 |5.23E+13|  3.56E-05|+/-4.60E-06|Jy|2005ApJ...635..853B|uncertainty|   5.731   microns   | Broad-band measurement|123707.21 +621408.1 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged new and previously published data
31|5.8 microns (IRAC)  | 32.7      |+/-3.9  |microJy             |5.23E+13|  3.27E-05|+/-3.90E-06|Jy|2009ApJ...699.1610H|uncertainty|     5.731 microns   | Broad-band measurement|12 37 07.20 +62 14 08.0 (J2000)| Flux in fixed aperture|                                        |From new raw data
32|PAH 6.2 (Spitzer)   | 1.41E-15  |+/-0.37E-15|erg/s/cm^2^         |4.84E+13|  1.41E+08|+/-3.70E+07|Jy-Hz|2009ApJ...699..667M|rms uncertainty|       6.2 microns   | Line measurement; flux integrated over line; lines measured in emission|12 37 07.21 +62 14 08.1 (J2000)| Flux integrated from map|                                        |From new raw data
33|PAH 7.7 (Spitzer)   | 3.53E-15  |+/-0.49E-15|erg/s/cm^2^         |3.89E+13|  3.53E+08|+/-4.90E+07|Jy-Hz|2009ApJ...699..667M|rms uncertainty|       7.7 microns   | Line measurement; flux integrated over line; lines measured in emission|12 37 07.21 +62 14 08.1 (J2000)| Flux integrated from map|                                        |From new raw data
34|8.0 microns (IRAC)  | 29.1      |+/-3.0  |microJy             |3.85E+13|  2.91E-05|+/-3.00E-06|Jy|2009ApJ...699.1610H|uncertainty|     7.782 microns   | Broad-band measurement|12 37 07.20 +62 14 08.0 (J2000)| Flux in fixed aperture|                                        |From new raw data
35|8.0 microns IRAC AB | 20.30     |+/-0.05 |mag                 |3.81E+13|  2.75E-05|+/-1.27E-06|Jy|2005ApJ...635..853B|uncertainty|   7.872   microns   | Broad-band measurement|123707.21 +621408.1 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged new and previously published data
36|PAH 8.6 (Spitzer)   | 0.83E-15  |+/-0.22E-15|erg/s/cm^2^         |3.49E+13|  8.30E+07|+/-2.20E+07|Jy-Hz|2009ApJ...699..667M|rms uncertainty|       8.6 microns   | Line measurement; flux integrated over line; lines measured in emission|12 37 07.21 +62 14 08.1 (J2000)| Flux integrated from map|                                        |From new raw data
37|16 microns (Spitzer)||<0.02      | milliJy            |1.87E+13||2.00E-05|Jy|2008ApJ...675.1171P|no uncertainty reported|        16 microns   | Broad-band measurement|12 37 07.19 +62 14 08.0 (J2000)| Flux integrated from map|                                        |Averaged from previously published data
38|24 microns (MIPS)   | 247.0     |+/-26.0 |microJy             |1.27E+13|  2.47E-04|+/-2.60E-05|Jy|2009ApJ...699.1610H|uncertainty|     23.68 microns   | Broad-band measurement|123707.21 +621408.1 (J2000)| Flux in fixed aperture|                                        |From new raw data
39|24 microns (MIPS)   | 255.0     |+/-9.0 |microJy              |1.27E+13|  2.55E-04|+/-9.0E-06|Jy|2009ApJ...699.1610H|uncertainty|     23.68 microns   | Broad-band measurement|123707.21 +621408.1 (J2000)| Flux in fixed aperture|                                        |From new raw data
40|24 microns (Spitzer)| 235       |+/-8    |microJy             |1.27E+13|  2.35E-04|+/-8.00E-06|Jy|2011ApJ...726...93R|uncertainty|     23.68 microns   | Broad-band measurement|12 37 07.21 +62 14 08.1 (J2000)| Not reported in paper|                                        |Averaged from previously published data
41|70 microns (Spitzer)||<3.5       | milliJy            |4.20E+12||3.50E-03|Jy|2008ApJ...675.1171P|no uncertainty reported|     71.42 microns   | Broad-band measurement|12 37 07.19 +62 14 08.0 (J2000)| Flux integrated from map|                                        |Averaged from previously published data
42|70 microns (MIPS)   ||<1.6       |microJy             |4.20E+12||1.60E-06|Jy|2009ApJ...699.1610H|3 sigma|     71.42 microns   | Broad-band measurement|123707.21 +621408.1 (J2000)| Flux in fixed aperture|                                        |From new raw data
43|70 microns (PACS)  |           |<2.0    |mJy                 |4.283E+12|         |2.0E-03|Jy|2004MNRAS.354..779G|3sigma uncertainty|      1200 microns   | Broad-band measurement|16 36 55.9 +40 59 12 (J2000)| Flux integrated from map|S/N = 3.66                              |From new raw data
44|100 microns (PACS) | 1.1       |+/-0.3  |microJy             |2.998e+12| 1.1E-03 |+/-0.3E-03 |Jy|2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
45|160 microns (PACS) | 6.4       |+/-1.3  |microJy             |1.874e+12| 6.4E-03 |+/-1.3E-03 |Jy|2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
46|250 microns (SPIRE)| 23.9      |+/-4.6  |mJy                 |1.199e+12| 23.9E-03 |+/-4.6e-03 |Jy|2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
47|350 microns (SPIRE)| 28.3      |+/-6.4  |mJy                 |8.565E+11| 28.3E-03 |+/-6.4E-03|Jy|2004MNRAS.354..779G|3sigma uncertainty|      1200 microns   | Broad-band measurement|16 36 55.9 +40 59 12 (J2000)| Flux integrated from map|S/N = 3.66                              |From new raw data
48|500 microns (SPIRE)| 23.8      |+/-4.0  |mJy                 |5.996E+11| 23.8E-03 |+/-4.0E-03|Jy|2004MNRAS.354..779G|3sigma uncertainty|      1200 microns   | Broad-band measurement|16 36 55.9 +40 59 12 (J2000)| Flux integrated from map|S/N = 3.66                              |From new raw data
49|850 microns (SCUBA) | 10.7     |+/-2.7  |milliJy             |3.53E+11|  1.07E-02|+/-2.70E-03|Jy|2005MNRAS.358..149P|uncertainty|     850   microns   | Broad-band measurement|12 37 07.7 +62 14 11 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
50|850 microns (SCUBA) | 8.0      |+/-3.1  |milliJy             |3.53E+11|  8.0E-03|+/-3.10E-03|Jy|2005MNRAS.358..149P|uncertainty|     850   microns   | Broad-band measurement|12 37 07.7 +62 14 11 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
51|850 microns (SCUBA) | 4.7      |+/-1.5  |milliJy             |3.53E+11|  4.70E-03|+/-1.50E-03|Jy|2005ApJ...622..772C|uncertainty|     850   microns   | Broad-band measurement|123707.21 +621408.1 (J2000)| Flux integrated from map|                                        |From new raw data
52|1160 microns (Penner)|         |<1.6    |mJy                 |2.58442E+11|       |1.6E-03|Jy|2004MNRAS.354..779G|3sigma uncertainty|      1200 microns   | Broad-band measurement|16 36 55.9 +40 59 12 (J2000)| Flux integrated from map|S/N = 3.66                              |From new raw data
52|1.3 mm (PdBI)       ||<1.4       |milliJy             |2.31E+11||1.40E-03|Jy|2006ApJ...640..228T|no uncertainty reported|     1.3   mm        | Broad-band measurement|| Flux integrated from map|                                        |From new raw data
54|8.5 GHz             | 16.20     ||microJy             |8.50E+09|  1.62E-05||Jy|1998AJ....116.1039R|no uncertainty reported|8.5        GHz       | Broad-band measurement; broad-band flux derived by integration over spectrum; synthetic band|123707.204 +621408.17 (J2000)| Flux integrated from map; Pointing and beam filling|                                        |From new raw data; Corrected for contaminating sources
55|8.5 GHz             | 15.90     ||microJy             |8.50E+09|  1.59E-05||Jy|1998AJ....116.1039R|no uncertainty reported|8.5        GHz       | Broad-band measurement; peak value reported; synthetic band|123707.204 +621408.17 (J2000)| Flux integrated from map; Pointing and beam filling|                                        |From new raw data; Corrected for contaminating sources
56|1.4 GHz (VLA)       | 28.3      |+/-4.2  |microJy             |1.40E+09|  2.83E-05|+/-4.20E-06|Jy|2010ApJS..188..178M|uncertainty|       1.4 GHz       | Broad-band measurement|12 37 07.18 +62 14 08.2 (J2000)| Total flux; Beam filling or dilution corrected|Major=0.0"; Minor=0.0"; PA=0 deg        |From new raw data
57|1.4 GHz             | 45.3      |+/-7.9  |microJy             |1.40E+09|  4.53E-05|+/-7.90E-06|Jy|2000ApJ...533..611R|1 sigma|1.4        GHz       | Broad-band measurement; broad-band flux derived by integration over spectrum; synthetic band|123707.208 +621408.08 (J2000)| Flux integrated from map; Pointing and beam filling|                                        |From new raw data; Corrected for contaminating sources
58|1.4 GHz (VLA)       | 45        ||microJy             |1.40E+09|  4.50E-05||Jy|2005MNRAS.358.1159M|no uncertainty reported|     1.4   GHz       | Broad-band measurement|12 37 07.2209 +62 14 08.208 (J2000)| Flux integrated from map|                                        |From new raw data
59|1.4 GHz (VLA)       | 39.      |+/-8.  | microJy            |1.40E+09|  39.E-06|+/-8.E-06|Jy|2007MNRAS.380..199I|rms uncertainty|       1.4 GHz       | Broad-band measurement|10 52 28.995 +57 22 22.42 (J2000)| Flux integrated from map|                                        |From reprocessed raw data
