
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-04-04T09:09:18PDT



Photometric Data for MM J163706+4053

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|[O II] 3727 (SUBARU)| 1.0E-16   |+/-0.3E-16|ergs cm^-2^ s^-1^   |8.04E+14|  1.24E-08|+/-3.73E-09|Jy|2006ApJ...651..713T|uncertainty|    3727   A         | Line measurement; flux integrated over line; lines measured in emission| | Flux integrated from map|                                        |From new raw data
2|H{beta} (SUBARU)    | 0.6E-16   |+/-0.3E-16|ergs cm^-2^ s^-1^   |6.17E+14|  9.72E-09|+/-4.86E-09|Jy|2006ApJ...651..713T|uncertainty|    4861   A         | Line measurement; flux integrated over line; lines measured in emission| | Flux integrated from map|                                        |From new raw data
3|[O III] 4959 SUBARU | 1.9E-16   |+/-0.6E-16|ergs cm^-2^ s^-1^   |6.05E+14|  3.14E-08|+/-9.92E-09|Jy|2006ApJ...651..713T|uncertainty|    4959   A         | Line measurement; flux integrated over line; lines measured in emission| | Flux integrated from map|                                        |From new raw data
4|[O III] 5007 SUBARU | 5.7E-16   |+/-0.6E-16|ergs cm^-2^ s^-1^   |5.99E+14|  9.52E-08|+/-1.00E-08|Jy|2006ApJ...651..713T|uncertainty|    5007   A         | Line measurement; flux integrated over line; lines measured in emission| | Flux integrated from map|                                        |From new raw data
5|H{alpha} (SUBARU)   | 7.4E-16   |+/-1.4E-16|ergs cm^-2^ s^-1^   |4.57E+14|  1.62E-07|+/-3.06E-08|Jy|2006ApJ...651..713T|uncertainty|    6563   A         | Line measurement; flux integrated over line; lines measured in emission| | Flux integrated from map|                                        |From new raw data
6|H{alpha} (Keck)     | 4.7E-19   |+/-0.6E-19| W/m^2^             |4.57E+14|  1.03E-07|+/-1.31E-08|Jy|2004ApJ...617...64S|uncertainty|      6563 A         | Line measurement; flux integrated over line; lines measured in emission|163706.51 +405313.8 (J2000)| Flux integrated from map|                                        |From new raw data
7|H{alpha} (Keck)     | 2.7E-19   |+/-0.8E-19| W/m^2^             |4.57E+14|  5.91E-08|+/-1.75E-08|Jy|2004ApJ...617...64S|uncertainty|      6563 A         | Line measurement; flux integrated over line; lines measured in emission|163706.51 +405313.8 (J2000)| Flux integrated from map|Broad-line component                    |From new raw data
6|F775W (HST/NICMOS)  | 24.40    |+/-0.06| mag                |3.93E+14| 6.30958e-07|+/-3.4868007e-08|Jy|2007A&A...470..467C|internal error|       1.6 microns   | Broad-band measurement| | From fitting to map|                                        |From new raw data
8|I (Cousins)         | 23.18     |+/-0.13 |mag                 |3.79E+14|  1.36E-06|+/-1.73E-07|Jy|2004ApJ...616...71S|1 sigma|    7900   A         | Broad-band measurement| | Flux in fixed aperture|4" aper; phot contam by near neighbor   |Averaged new and previously published data
3|HST F110W            | 23.66     |+/-0.07 |mag             |2.67195e+14|1.24738e-06|+/-8.0421731e-08|Jy |2011ApJ...728L...4H|uncertainty|     3.550 microns   | Broad-band measurement|09 03 11.6 +00 39 06 (J2000)| Flux in fixed aperture|                                        |From new raw data
6|F160W (HST/NICMOS)  | 21.93    |+/-0.01| mag                |1.87E+14| 6.13761e-06|+/-5.6529522e-08|Jy|2007A&A...470..467C|internal error|       1.6 microns   | Broad-band measurement| | From fitting to map|                                        |From new raw data
9|K_s_ (2MASS)        | 19.16     |+/-0.06 |mag                 |1.38E+14|  1.44E-05|+/-8.21E-07|Jy|2004ApJ...616...71S|1 sigma|    2.17   microns   | Broad-band measurement| | Flux in fixed aperture|4" aper; phot contam by near neighbor   |Averaged new and previously published data
10|4.5 microns (IRAC)  | 32.4      |+/-3.3  |microJy             |6.67E+13|  3.24E-05|+/-3.30E-06|Jy|2009ApJ...699.1610H|uncertainty|     4.493 microns   | Broad-band measurement|16 37 06.47 +40 53 14.2 (J2000)| Flux in fixed aperture|                                        |From new raw data
11|7.7 microns (IRS)   | 0.519     | |milliJy             |3.89E+13|  5.19E-04| |Jy|2007ApJ...660.1060V|no uncertainty reported|     7.7   microns   | Line measurement; flux integrated over line; lines measured in emission|16 37 06.60 +40 53 14.0 (J2000)| Flux integrated from map|                                        |From new raw data
12|7.7 microns (IRS)   | 0.242     | |milliJy             |3.89E+13|  2.42E-04| |Jy|2007ApJ...660.1060V|no uncertainty reported|     7.7   microns   | Broad-band measurement|16 37 06.60 +40 53 14.0 (J2000)| Flux integrated from map|                                        |From new raw data
13|8.0 microns (IRAC)  | 63.8      |+/-6.5  |microJy             |3.85E+13|  6.38E-05|+/-6.50E-06|Jy|2009ApJ...699.1610H|uncertainty|     7.782 microns   | Broad-band measurement|16 37 06.47 +40 53 14.2 (J2000)| Flux in fixed aperture|                                        |From new raw data
14|24 microns (MIPS)   | 0.41      |+/-10  %|milliJy             |1.27E+13|  4.10E-04|+/-4.10E-05|Jy|2009A&A...502..541E|uncertainty|     23.68 microns   | Broad-band measurement| | Flux in fixed aperture|                                        |From reprocessed raw data
15|24 microns (MIPS)   | 375.0     |+/-60.0 |microJy             |1.27E+13|  3.75E-04|+/-6.00E-05|Jy|2009ApJ...699.1610H|uncertainty|     23.68 microns   | Broad-band measurement|163706.51 +405313.8 (J2000)| Flux in fixed aperture|                                        |From new raw data
16|70 microns (MIPS)   | |<5.1       |milliJy             |4.20E+12| |5.10E-03|Jy|2009A&A...502..541E|3 sigma|     71.42 microns   | Broad-band measurement| | Flux in fixed aperture|                                        |From reprocessed raw data
17|70 microns (MIPS)   | |<9.5       |milliJy             |4.20E+12| |9.50E-03|Jy|2009ApJ...699.1610H|3 sigma|     71.42 microns   | Broad-band measurement|163706.51 +405313.8 (J2000)| Flux in fixed aperture|                                        |From new raw data
18|160 microns (MIPS)  | |<17        |milliJy             |1.92E+12| |1.70E-02|Jy|2009A&A...502..541E|3 sigma|     155.9 microns   | Broad-band measurement| | Flux in fixed aperture|                                        |From reprocessed raw data
19|350 microns (SHARC2)| 36.1      |+/-7.7  |milliJy             |8.57E+11|  3.61E-02|+/-7.70E-03|Jy|2006ApJ...650..592K|uncertainty|     350   microns   | Broad-band measurement| | Total flux|                                        |From new raw data
20|850 microns (SCUBA) | 11.2      |+/-2.9  |milliJy             |3.53E+11|  1.12E-02|+/-2.90E-03|Jy|2005ApJ...622..772C|uncertainty|     850   microns   | Broad-band measurement|163706.51 +405313.8 (J2000)| Flux integrated from map|                                        |From new raw data
21|CO(3-2) line (IRAM) | 1.0       |+/-0.2  |Jy km s^-1^         |3.46E+11|  2.92E-07|+/-5.84E-08|Jy|2005MNRAS.359.1165G|uncertainty|   2.380             | Line measurement; flux integrated over line; lines measured in emission|16 37 06.50 +40 53 13.8 (J2000)| Flux integrated from map|                                        |From new raw data
22|1200 microns (MAMBO)| 4.2       |+/-1.1  | milliJy            |2.50E+11|  4.20E-03|+/-1.10E-03|Jy|2004MNRAS.354..779G|uncertainty|      1200 microns   | Broad-band measurement|16 37 06.7 +40 53 15 (J2000)| Flux integrated from map|S/N = 3.81                              |From new raw data
