
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-07-10T13:42:15PDT



Photometric Data for SPT-SJ214654-5507.8

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
6|24 microns (MIPS)   | 150.0     |+/-15.0  |microJy             |1.27E+13|  150.0E-06|+/-15.0E-06|Jy|2011AJ....141....1T|rms uncertainty|     23.68 microns   | Broad-band measurement|189.110626 62.143169 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
5|250 microns (SPIRE)| 19.0      |+/-3.4 |mJy             |1.199e+12| 19.0E-03|+/-3.4e-03 |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
6|350 microns (SPIRE)| 18.7      |+/-3.7  |mJy             |8.565e+11|18.7E-03 |+/-3.7e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
8|500 microns (SPIRE) |      |<10.4 |mJy             |5.996e+11||10.4E-03 |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
