
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-07-13T02:04:37PDT



Photometric Data for GOODS J123712.04+621212.3

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|4.0-8 keV (Chandra) ||<0.45E-15  |ergs cm^-2^ s^-1^   |1.45E+18||3.10E-11|Jy|2003AJ....126..539A|3 sigma|       6   keV       | Broad-band measurement|12 37 12.09 +62 12 11.3 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
2|4-8 keV (Chandra)   ||<0.46E-15  |erg cm^-2^ s^-1^    |1.45E+18||3.17E-11|Jy|2001AJ....122.2810B|no uncertainty reported|       6   keV       | Broad-band measurement|12 37 12.11 +62 12 11.3 (J2000)| Flux in fixed aperture|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
3|2-8 keV (Chandra)   | 0.27E-15  |+/-4   %|erg cm^-2^ s^-1^    |1.21E+18|  2.23E-11|+/-8.93E-13|Jy|2001AJ....122.2810B|estimated error|       5   keV       | Broad-band measurement|12 37 12.11 +62 12 11.3 (J2000)| Flux in fixed aperture|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
4|2.0-8 keV (Chandra) | 0.37E-15  ||ergs cm^-2^ s^-1^   |1.21E+18|  3.06E-11||Jy|2003AJ....126..539A|no uncertainty reported|       5   keV       | Broad-band measurement|12 37 12.09 +62 12 11.3 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
5|0.5-8 keV (Chandra) | 0.19E-15  |+/-4   %|erg cm^-2^ s^-1^    |1.03E+18|  1.84E-11|+/-7.38E-13|Jy|2001AJ....122.2810B|estimated error|    4.25   keV       | Broad-band measurement|12 37 12.11 +62 12 11.3 (J2000)| Flux in fixed aperture|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
6|0.5-8 keV (Chandra) | 0.38E-15  ||ergs cm^-2^ s^-1^   |1.03E+18|  3.70E-11||Jy|2003AJ....126..539A|no uncertainty reported|    4.25   keV       | Broad-band measurement|12 37 12.09 +62 12 11.3 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
7|2.0-4 keV (Chandra) ||<0.12E-15  |ergs cm^-2^ s^-1^   |7.25E+17||1.65E-11|Jy|2003AJ....126..539A|3 sigma|       3   keV       | Broad-band measurement|12 37 12.09 +62 12 11.3 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
8|1.0-2 keV (Chandra) | 0.02E-15  ||ergs cm^-2^ s^-1^   |3.63E+17|  5.51E-12||Jy|2003AJ....126..539A|no uncertainty reported|     1.5   keV       | Broad-band measurement|12 37 12.09 +62 12 11.3 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
9|0.5-2 keV (Chandra) | 0.03E-15  ||ergs cm^-2^ s^-1^   |3.02E+17|  9.92E-12||Jy|2003AJ....126..539A|no uncertainty reported|    1.25   keV       | Broad-band measurement|12 37 12.09 +62 12 11.3 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
10|0.5-2 keV (Chandra) ||<0.05E-15  |erg cm^-2^ s^-1^    |3.02E+17||1.66E-11|Jy|2001AJ....122.2810B|no uncertainty reported|    1.25   keV       | Broad-band measurement|12 37 12.11 +62 12 11.3 (J2000)| Flux in fixed aperture|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
11|0.5-1 keV (Chandra) ||<0.04E-15  |ergs cm^-2^ s^-1^   |1.81E+17||2.21E-11|Jy|2003AJ....126..539A|3 sigma|    0.75   keV       | Broad-band measurement|12 37 12.09 +62 12 11.3 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
12|U (KPNO/MOSAIC) AB  ||>27.8      |mag                 |8.44E+14||2.75E-08|Jy|2005ApJ...635..853B|2.5 sigma|    3552   A         | Broad-band measurement|123712.05 +621212.3 (J2000)| Flux in fixed aperture|3" aperture                             |Averaged new and previously published data
13|F435W (HST) AB      | 29.292    ||mag                 |6.98E+14|  6.97E-09||Jy|2010A&A...522A..11R|no uncertainty reported|      4297 A         | Broad-band measurement|189.300284 62.203440 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
14|B (Subaru) AB       ||>27.6      |mag                 |6.81E+14||3.31E-08|Jy|2005ApJ...635..853B|2.5 sigma|    4400   A         | Broad-band measurement|123712.05 +621212.3 (J2000)| Flux in fixed aperture|3" aperture                             |Averaged new and previously published data
15|V (Subaru) AB       ||>27.6      |mag                 |5.42E+14||3.31E-08|Jy|2005ApJ...635..853B|2.5 sigma|    5530   A         | Broad-band measurement|123712.05 +621212.3 (J2000)| Flux in fixed aperture|3" aperture                             |Averaged new and previously published data
16|F606W (HST) AB      | 28.546    ||mag                 |5.08E+14|  1.39E-08||Jy|2010A&A...522A..11R|no uncertainty reported|      5907 A         | Broad-band measurement|189.300284 62.203440 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
17|R (Subaru) AB       ||>27.4      |mag                 |4.68E+14||3.98E-08|Jy|2005ApJ...635..853B|2.5 sigma|    6400   A         | Broad-band measurement|123712.05 +621212.3 (J2000)| Flux in fixed aperture|3" aperture                             |Averaged new and previously published data
18|F775W (HST) AB      | 27.613    ||mag                 |3.86E+14|  3.27E-08||Jy|2010A&A...522A..11R|no uncertainty reported|      7764 A         | Broad-band measurement|189.300284 62.203440 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
19|I (Subaru) AB       ||>26.4      |mag                 |3.79E+14||1.00E-07|Jy|2005ApJ...635..853B|2.5 sigma|    7900   A         | Broad-band measurement|123712.05 +621212.3 (J2000)| Flux in fixed aperture|3" aperture                             |Averaged new and previously published data
20|I (Cousins)         | 25.71     |+/-0.33 |mag                 |3.79E+14|  1.33E-07|+/-4.71E-08|Jy|2004ApJ...616...71S|1 sigma|    7900   A         | Broad-band measurement|| Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
21|z' (Subaru) AB      ||>26.2      |mag                 |3.30E+14||1.20E-07|Jy|2005ApJ...635..853B|2.5 sigma|    9097   A         | Broad-band measurement|123712.05 +621212.3 (J2000)| Flux in fixed aperture|3" aperture                             |Averaged new and previously published data
22|F850LP (HST) AB     | 27.172    ||mag                 |3.17E+14|  4.91E-08||Jy|2010A&A...522A..11R|no uncertainty reported|      9445 A         | Broad-band measurement|189.300284 62.203440 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
23|J (2MASS)           ||>22.50     |mag                 |2.40E+14||1.59E-06|Jy|2004ApJ...616...71S|3sigma uncertainty|    1.25   microns   | Broad-band measurement|| Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
24|J (Hale/WIRC) AB    ||>24.0      |mag                 |2.40E+14||9.12E-07|Jy|2005ApJ...635..853B|2.5 sigma|   1.250   microns   | Broad-band measurement|123712.05 +621212.3 (J2000)| Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
25|F160W (HST) AB      | 23.21     |+/-0.13 |mag                 |1.87E+14|  1.89E-06|+/-2.26E-07|Jy|2011MNRAS.413...80C|uncertainty|      1.60 microns   | Broad-band measurement|189.300201 62.203414 (J2000)| Total flux|                                        |From new raw data
26|HK' (UH:2.2m) AB    | 21.945    ||mag                 |1.59E+14|  6.05E-06||Jy|2010A&A...522A..11R|no uncertainty reported|      1.89 microns   | Broad-band measurement|189.300284 62.203440 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
27|K_s (Hale/WIRC) AB  | 23.02     |+/-0.30 |mag                 |1.39E+14|  2.25E-06|+/-6.22E-07|Jy|2005ApJ...635..853B|uncertainty|   2.150   microns   | Broad-band measurement|123712.05 +621212.3 (J2000)| Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
28|K_s (Hale/WIRC) AB  | 22.47     ||mag                 |1.39E+14|  3.73E-06||Jy|2005ApJ...633..748R|no uncertainty reported|   2.150   microns   | Broad-band measurement|12 37 12.05 +62 12 12.3 (J2000)| Flux in fixed aperture|                                        |From new raw data
29|K_s (Subaru)        | 20.728    ||mag                 |1.39E+14|  3.46E-06||Jy|2010A&A...522A..11R|no uncertainty reported|      2.15 microns   | Broad-band measurement|189.300284 62.203440 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
30|K_s (2MASS)         | 20.76     |+/-0.32 |mag                 |1.38E+14|  3.31E-06|+/-1.14E-06|Jy|2004ApJ...616...71S|1 sigma|    2.17   microns   | Broad-band measurement|| Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
31|3.6 microns (IRAC)  | 11.1      |+/-1.3  |microJy             |8.44E+13|  1.11E-05|+/-1.30E-06|Jy|2009ApJ...699.1610H|uncertainty|     3.550 microns   | Broad-band measurement|12 37 12.05 +62 12 11.9 (J2000)| Flux in fixed aperture|                                        |From new raw data
32|3.6 microns (IRAC)  | 10.584    ||microJy             |8.44E+13|  1.06E-05||Jy|2010A&A...522A..11R|no uncertainty reported|     3.550 microns   | Broad-band measurement|189.300284 62.203440 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
33|4.5 microns IRAC AB | 29.95     |+/-0.07 |mag                 |6.67E+13|  3.80E-09|+/-2.45E-10|Jy|2005ApJ...635..853B|uncertainty|   4.493   microns   | Broad-band measurement|123712.05 +621212.3 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged new and previously published data
34|4.5 microns (IRAC)  | 15.2      |+/-1.5  |microJy             |6.67E+13|  1.52E-05|+/-1.50E-06|Jy|2009ApJ...699.1610H|uncertainty|     4.493 microns   | Broad-band measurement|12 37 12.05 +62 12 11.9 (J2000)| Flux in fixed aperture|                                        |From new raw data
35|4.5 microns (IRAC)  | 14.332    ||microJy             |6.67E+13|  1.06E-05||Jy|2010A&A...522A..11R|no uncertainty reported|     4.493 microns   | Broad-band measurement|189.300284 62.203440 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
36|5.8 microns IRAC AB | 20.62     |+/-0.13 |mag                 |5.23E+13|  2.05E-05|+/-2.46E-06|Jy|2005ApJ...635..853B|uncertainty|   5.731   microns   | Broad-band measurement|123712.05 +621212.3 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged new and previously published data
37|5.8 microns (IRAC)  | 21.3      |+/-2.2  |microJy             |5.23E+13|  2.13E-05|+/-2.20E-06|Jy|2009ApJ...699.1610H|uncertainty|     5.731 microns   | Broad-band measurement|12 37 12.05 +62 12 11.9 (J2000)| Flux in fixed aperture|                                        |From new raw data
38|5.8 microns (IRAC)  | 21.049    ||microJy             |5.23E+13|  2.11E-05||Jy|2010A&A...522A..11R|no uncertainty reported|     5.731 microns   | Broad-band measurement|189.300284 62.203440 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
39|8.0 microns (IRAC)  | 24.2      |+/-2.5  |microJy             |3.85E+13|  2.42E-05|+/-2.50E-06|Jy|2009ApJ...699.1610H|uncertainty|     7.782 microns   | Broad-band measurement|12 37 12.05 +62 12 11.9 (J2000)| Flux in fixed aperture|                                        |From new raw data
40|8.0 microns IRAC AB | 20.58     |+/-0.05 |mag                 |3.81E+13|  2.13E-05|+/-9.80E-07|Jy|2005ApJ...635..853B|uncertainty|   7.872   microns   | Broad-band measurement|123712.05 +621212.3 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged new and previously published data
41|8.0 microns (IRAC)  | 20.979    ||microJy             |3.81E+13|  2.10E-05||Jy|2010A&A...522A..11R|no uncertainty reported|     7.872 microns   | Broad-band measurement|189.300284 62.203440 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
42|24 microns (MIPS)   | 30.0      |+/-8.6  |microJy             |1.27E+13|  3.00E-05|+/-8.60E-06|Jy|2009ApJ...699.1610H|uncertainty|     23.68 microns   | Broad-band measurement|123712.05 +621212.3 (J2000)| Flux in fixed aperture|                                        |From new raw data
43|24 microns (MIPS)   ||<80.0      |microJy             |1.27E+13||8.00E-05|Jy|2007ApJ...660..167D|no uncertainty reported|   23.68   microns   | Broad-band measurement|12 37 12.07 +62 12 11.61 (J2000)| Flux in fixed aperture|                                        |From new raw data
44|24 microns (MIPS)   | 48.774    ||microJy             |1.27E+13|  4.88E-05||Jy|2010A&A...522A..11R|no uncertainty reported|     23.68 microns   | Broad-band measurement|189.300284 62.203440 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
45|24 microns (MIPS)   | 51.3      |+/-2.7  |microJy             |1.27E+13|  5.13E-05|+/-2.70E-06|Jy|2011A&A...528A..35M|uncertainty|     23.68 microns   | Broad-band measurement|12 37 12.05 +62 12 11.91 (J2000)| Flux integrated from map|                                        |From new raw data
46|70 microns (MIPS)   ||<1.5       |microJy             |4.20E+12||1.50E-06|Jy|2009ApJ...699.1610H|3 sigma|     71.42 microns   | Broad-band measurement|123712.05 +621212.3 (J2000)| Flux in fixed aperture|                                        |From new raw data
47|70 microns (MIPS)   ||<2.1       |milliJy             |4.20E+12||2.10E-03|Jy|2011A&A...528A..35M|no uncertainty reported|     71.42 microns   | Broad-band measurement|12 37 12.05 +62 12 11.91 (J2000)| Flux integrated from map|                                        |From new raw data
48|850 microns (SCUBA) | 8.0       |+/-1.8  |milliJy             |3.53E+11|  8.00E-03|+/-1.80E-03|Jy|2005ApJ...622..772C|uncertainty|     850   microns   | Broad-band measurement|123712.05 +621212.3 (J2000)| Flux integrated from map|                                        |From new raw data
1|850um (SCUBA)   | 8.0 |+/-1.8| mJy  | 3.529E11| 8.0E-3| 1.8E-3 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
49|340 GHz (SMA)       | 5.34      |+/-0.97 |milliJy             |3.40E+11|  5.34E-03|+/-9.70E-04|Jy|2011ApJ...726L..18W|uncertainty|       340 GHz       | Broad-band measurement|189.30002 62.20341 (J2000)| Flux integrated from map|Primary beam corrected                  |From new raw data
50|1.4 GHz (VLA)       | 31.7      |+/-4.3  |microJy             |1.40E+09|  3.17E-05|+/-4.30E-06|Jy|2010ApJS..188..178M|uncertainty|       1.4 GHz       | Broad-band measurement|12 37 12.04 +62 12 11.7 (J2000)| Total flux; Beam filling or dilution corrected|Major=0.5"; Minor=0.0"; PA=135 deg      |From new raw data
2|1.4GHz (VLA)    | 21.0|+/-4.0| uJy  | 1.4E9| 21.0E-6| 4.0E-6 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
