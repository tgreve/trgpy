
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-07-10T07:03:41PDT



Photometric Data for BRI 1335-0417

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|[CII] 157.74 (APEX) | 26.6      |+/-4.3  |Jy km/s             |1.90E+12|  3.12E+07|+/-5.04E+06|Jy-Hz|2010A&A...519L...1W|uncertainty|    157.74 microns   | Line measurement; flux integrated over line; lines measured in emission|13 38 03.38 -04 32 35.3 (J2000)| Total flux|                                        |From new raw data
2|350 microns (SHARC-II)        | 0.052     |+/-0.008|Jy                  |8.57E+11|  5.20E-02|+/-8.00E-03|Jy|1999CIT...T00R....B|1 sigma|350        microns   | Broad-band measurement|133527.6 -041721. (B1950)| Flux integrated from map|                                        |From new raw data
3|CI(2-1) (IRAM 30)   ||<0.8       |Jy km/s             |8.09E+11||3.99E+05|Jy-Hz|2011ApJ...730...18W|5 sigma|   809.344 GHz       | Line measurement; flux integrated over line; lines measured in emission|13 38 03.42 -04 32 34.1 (J2000)| Flux integrated from map|                                        |From new raw data
4|CI(1-0) (IRAM 30)   ||<2.2       |Jy km/s             |4.92E+11||6.68E+05|Jy-Hz|2011ApJ...730...18W|3 sigma|   492.161 GHz       | Line measurement; flux integrated over line; lines measured in emission|13 38 03.42 -04 32 34.1 (J2000)| Flux integrated from map|                                        |From new raw data
5|1.4 GHz (VLBI)      | 208       |+/-46   | microJy            |1.40E+09|  2.08E-04|+/-4.60E-05|Jy|2007AJ....134..694M|uncertainty|    1.4    GHz       | Broad-band measurement|| Total flux|                                        |From new raw data
