
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-06-14T16:43:48PDT



Photometric Data for PKS 1623+26:[SSP2004] BX0453

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|G (WHT)             | 23.86     ||mag                 |6.38E+14|  1.04E-06||Jy|2006ApJ...647..128E|no uncertainty reported|    0.47   microns   | Broad-band measurement|| Flux in fixed aperture|                                        |Averaged from previously published data
9|J (Hale/WIRC)       | 21.41     ||mag                 |2.40E+14|  4.26E-06||Jy|2006ApJ...646..107E|no uncertainty reported|    1.25   microns   | Broad-band measurement|16 25 50.84 +26 49 31.40 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data; derived from aflux in a different band and a color
10|K_s (Hale/WIRC)     | 19.76     ||mag                 |1.39E+14|  8.36E-06||Jy|2006ApJ...646..107E|no uncertainty reported|    2.15   microns   | Broad-band measurement|16 25 50.84 +26 49 31.40 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data
11|3.6 microns IRAC AB | 21.38     || mag                |8.44E+13|  1.02E-05||Jy|2007ApJ...669..929L|no uncertainty reported|     3.550 microns   | Broad-band measurement|16 25 50.854 +26 49 31.28 (J2000)| Flux integrated from map|                                        |From reprocessed raw data
12|4.5 microns IRAC AB | 21.37     || mag                |6.67E+13|  1.03E-05||Jy|2007ApJ...669..929L|no uncertainty reported|     4.493 microns   | Broad-band measurement|16 25 50.854 +26 49 31.28 (J2000)| Flux integrated from map|                                        |From reprocessed raw data
13|5.8 microns IRAC AB | 21.33     || mag                |5.23E+13|  1.07E-05||Jy|2007ApJ...669..929L|no uncertainty reported|     5.731 microns   | Broad-band measurement|16 25 50.854 +26 49 31.28 (J2000)| Flux integrated from map|                                        |From reprocessed raw data
14|8.0 microns IRAC AB | 21.92     || mag                |3.81E+13|  6.20E-06||Jy|2007ApJ...669..929L|no uncertainty reported|     7.872 microns   | Broad-band measurement|16 25 50.854 +26 49 31.28 (J2000)| Flux integrated from map|                                        |From reprocessed raw data
15|24 microns (MIPS)   | 195       || microJy            |1.27E+13|  1.95E-04||Jy|2007ApJ...669..929L|no uncertainty reported|     23.68 microns   | Broad-band measurement|16 25 50.854 +26 49 31.28 (J2000)| Flux integrated from map|                                        |From reprocessed raw data
