
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-07-08T08:37:11PDT



Photometric Data for 4C +05.19

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|0.5-8 keV (Chandra) | 13E-14    |+/-6E-14|ergs/cm^2^/s        |1.03E+18|  1.26E-08|+/-5.83E-09|Jy|2007ApJ...661...19P|uncertainty|    4.25   keV       | Broad-band measurement|| From fitting to map|Unabsorbed flux                         |From reprocessed raw data; NED frequency assigned tomid-point of band in keV
2|0.5-8 keV (Chandra) | 14E-14    |+/-4E-14|ergs/cm^2^/s        |1.03E+18|  1.36E-08|+/-3.88E-09|Jy|2007ApJ...661...19P|uncertainty|    4.25   keV       | Broad-band measurement|| From fitting to map|Unabsorbed flux                         |From reprocessed raw data; NED frequency assigned tomid-point of band in keV
3|0.5-8 keV (Chandra) | 12E-14    |+/-7E-14|ergs/cm^2^/s        |1.03E+18|  1.17E-08|+/-6.80E-09|Jy|2007ApJ...661...19P|uncertainty|    4.25   keV       | Broad-band measurement|| From fitting to map|Unabsorbed flux                         |From reprocessed raw data; NED frequency assigned tomid-point of band in keV
4|0.5-8 keV (Chandra) | 15E-14    |+/-6E-14|ergs/cm^2^/s        |1.03E+18|  1.46E-08|+/-5.83E-09|Jy|2007ApJ...661...19P|uncertainty|    4.25   keV       | Broad-band measurement|| From fitting to map|Unabsorbed flux                         |From reprocessed raw data; NED frequency assigned tomid-point of band in keV
5|0.5-8 keV (Chandra) | 14E-14    |+/-9E-14|ergs/cm^2^/s        |1.03E+18|  1.36E-08|+/-8.74E-09|Jy|2007ApJ...661...19P|uncertainty|    4.25   keV       | Broad-band measurement|| From fitting to map|Unabsorbed flux                         |From reprocessed raw data; NED frequency assigned tomid-point of band in keV
6|0.5-8 keV (Chandra) | 13E-14    |+/-3E-14|ergs/cm^2^/s        |1.03E+18|  1.26E-08|+/-2.91E-09|Jy|2007ApJ...661...19P|uncertainty|    4.25   keV       | Broad-band measurement|| From fitting to map|Unabsorbed flux                         |From reprocessed raw data; NED frequency assigned tomid-point of band in keV
7|0.5-8 keV (Chandra) | 16E-14    |+/-7E-14|ergs/cm^2^/s        |1.03E+18|  1.55E-08|+/-6.80E-09|Jy|2007ApJ...661...19P|uncertainty|    4.25   keV       | Broad-band measurement|| From fitting to map|Unabsorbed flux                         |From reprocessed raw data; NED frequency assigned tomid-point of band in keV
8|0.5-8 keV (Chandra) | 6.79E-13  |+/-0.33E-13|erg/cm^2^/s         |1.03E+18|  6.59E-08|+/-3.20E-09|Jy|2012ApJ...744..111P|uncertainty|      4.25 keV       | Broad-band measurement|| Total flux|                                        |From reprocessed raw data; Extinction-corrected for MilkyWay; NED frequency assigned to mid-point of band in keV
9|F555W (HST)         | 24.17     |+/-0.15 | mag                |5.54E+14|  8.01E-07|+/-1.11E-07|Jy|2008A&A...478...95Y|uncertainty|      5407 A         | Broad-band measurement|| Modelled datum|                                        |Averaged from previously published data
10|F814W (HST)         | 20.91     |+/-0.05 | mag                |3.78E+14|  1.08E-05|+/-4.96E-07|Jy|2008A&A...478...95Y|uncertainty|      7940 A         | Broad-band measurement|| Modelled datum|                                        |Averaged from previously published data
11|I (HST)             | 19.62     ||mag                 |3.68E+14|  3.42E-05||Jy|2011ApJ...738...96M|no uncertainty reported|     0.814 microns   | Broad-band measurement|| Not reported in paper|                                        |From reprocessed raw data
12|J_total (2MASS)     | 16.265    |+/-0.431|mag                 |2.40E+14|  4.97E-04|+/-2.42E-04|Jy|20032MASX.C.......:|1 sigma uncert.| 1.25      microns   | Broad-band measurement|041437.75 +053442.6 (J2000)| Total flux|                                        |From new raw data
13|J_14arcsec (2MASS)  | 16.265    |+/-0.431|mag                 |2.40E+14|  4.97E-04|+/-2.42E-04|Jy|20032MASX.C.......:|1 sigma uncert.| 1.25      microns   | Broad-band measurement|041437.75 +053442.6 (J2000)| Flux in fixed aperture|14.0 x 14.0 arcsec aperture.            |From new raw data
14|F160W (HST/NIC2)    | 18.63     ||mag                 |1.87E+14|  3.83E-05||Jy|2006ApJ...649..616P|no uncertainty reported|   1.606   microns   | Broad-band measurement|04 14 37.73 +05 34 44.3 (J2000)| From fitting to map|Quasar mag; extinction = 0.18           |From new raw data; Extinction-corrected for Milky Way
15|F160W (HST/NIC2)    | 20.78     |+/-0.3  |mag                 |1.87E+14|  5.28E-06|+/-4.31E-06|Jy|2006ApJ...649..616P|typical accuracy|   1.606   microns   | Broad-band measurement|04 14 37.73 +05 34 44.3 (J2000)| From fitting to map|Host mag; extinction = 0.18             |From new raw data; Extinction-corrected for Milky Way
16|F160W (HST)         | 17.54     |+/-0.14 | mag                |1.87E+14|  1.01E-04|+/-1.30E-05|Jy|2008A&A...478...95Y|uncertainty|     1.603 microns   | Broad-band measurement|| Modelled datum|                                        |Averaged from previously published data
17|H_total (2MASS)     | 14.158    |+/-0.103|mag                 |1.82E+14|  2.22E-03|+/-2.21E-04|Jy|20032MASX.C.......:|1 sigma uncert.| 1.65      microns   | Broad-band measurement|041437.75 +053442.6 (J2000)| Total flux|                                        |From new raw data
18|H_14arcsec (2MASS)  | 13.953    |+/-0.120|mag                 |1.82E+14|  2.69E-03|+/-3.14E-04|Jy|20032MASX.C.......:|1 sigma uncert.| 1.65      microns   | Broad-band measurement|041437.75 +053442.6 (J2000)| Flux in fixed aperture|14.0 x 14.0 arcsec aperture.            |From new raw data
19|H_K20 (2MASS)       | 14.158    |+/-0.103|mag                 |1.82E+14|  2.22E-03|+/-2.21E-04|Jy|20032MASX.C.......:|1 sigma uncert.| 1.65      microns   | Broad-band measurement|041437.75 +053442.6 (J2000)| Flux integrated from map|  10.0 x   10.0 arcsec integration area.|From new raw data
20|K_s_14arcsec (2MASS)| 13.628    |+/-0.159|mag                 |1.38E+14|  2.36E-03|+/-3.72E-04|Jy|20032MASX.C.......:|1 sigma uncert.| 2.17      microns   | Broad-band measurement|041437.75 +053442.6 (J2000)| Flux in fixed aperture|14.0 x 14.0 arcsec aperture.            |From new raw data
21|K_s                 | 13.715    |+/-0.123|mag                 |1.38E+14|  2.18E-03|+/-2.61E-04|Jy|20032MASX.C.......:|1 sigma uncert.| 2.17      cm        | Broad-band measurement|041437.75 +053442.6 (J2000)| Flux in fixed aperture|                                        |From new raw data
22|K_s                 | 13.715    |+/-0.123|mag                 |1.38E+14|  2.18E-03|+/-2.61E-04|Jy|20032MASX.C.......:|1 sigma uncert.| 2.17      cm        | Broad-band measurement|041437.75 +053442.6 (J2000)| Flux in fixed aperture|  10.0 x   10.0 arcsec integration area.|From new raw data
23|117 GHz             | 95.413    |+/-0.018 |Jy                  |1.17E+11| 95.413|+/-0.018|Jy|1973AJ.....78..828K|uncertainty|    10.7   GHz       | Broad-band measurement|| Total flux|                                        |From new raw data
23|10.7 GHz (NRAO)     | 0.38      |+/-0.02 |Jy                  |1.07E+10|  3.80E-01|+/-2.00E-02|Jy|1973AJ.....78..828K|uncertainty|    10.7   GHz       | Broad-band measurement|| Total flux|                                        |From new raw data
24|8.6 GHz (ATCA)      | 0.34      || Jy                 |8.60E+09|  3.40E-01||Jy|2003PASJ...55..351T|no uncertainty reported|       8.6 GHz       | Broad-band measurement|| Flux integrated from map|                                        |From new raw data
25|6.11 GHz (Arecibo)  | 0.71      |+/-0.02 |Jy                  |6.11E+09|  7.10E-01|+/-2.00E-02|Jy|2011A&A...529A.150C|uncertainty|      6.11 GHz       | Broad-band measurement|| Flux integrated from map|                                        |From new raw data
26|5000 MHz            | 0.710     ||Jy                  |5.00E+09|  7.10E-01||Jy|1990PKS90.C...0000W|no uncertainty reported|    5000   MHz       | Broad-band measurement|04 11 58.2 +05 27 13 (B1950)| Integrated from scans|                                        |Homogenized from new and previously published data
27|5 GHz (VLBA)        | 1.1       || Jy                 |5.00E+09|  1.10E+00||Jy|2004ApJ...616..110H|no uncertainty reported|         5 GHz       | Broad-band measurement|| Total flux|                                        |From new raw data
28|5 GHz (VLBI)        | 0.09      || Jy                 |5.00E+09|  9.00E-02||Jy|2008ApJS..175..314D|no uncertainty reported|         5 GHz       | Broad-band measurement|| Flux integrated from map|Core flux                               |Averaged new and previously published data
29|4.85 GHz            | 1110      |+/-154  |milliJy             |4.85E+09|  1.11E+00|+/-1.54E-01|Jy|1991ApJS...75.1011G|rms noise|4.85       GHz       | Broad-band measurement|041158.6 +052716 (B1950)| Modelled datum|                                        |From new raw data; Corrected for contaminating sources
30|4.85 GHz            | 959       |+/-51   |milliJy             |4.85E+09|  9.59E-01|+/-5.10E-02|Jy|1995ApJS...97..347G|rms noise|4.85       GHz       | Broad-band measurement|041437.4 +053438 (J2000)| Modelled datum|                                        |From new raw data; Corrected for contaminating sources
31|4.85 GHz            | 1119      |+/-15  %|milliJy             |4.85E+09|  1.12E+00|+/-1.68E-01|Jy|1991ApJS...75....1B|uncertainty|4.85       GHz       | Broad-band measurement|041158.7 +052718 (B1950)| Peak flux|                                        |From new raw data; Corrected for contaminating sources
32|4.8 GHz (ATCA)      | 0.68      || Jy                 |4.80E+09|  6.80E-01||Jy|2003PASJ...55..351T|no uncertainty reported|       4.8 GHz       | Broad-band measurement|| Flux integrated from map|                                        |From new raw data
33|4775 MHz (NRAO)     | 741       ||milliJy             |4.78E+09|  7.41E-01||Jy|1986ApJS...61....1B|no uncertainty reported|    4775   MHz       | Broad-band measurement|04 14 39.5 +05 34 35 (J2000)| Flux integrated from map|S/N = 41.0                              |From new raw data
34|2700 MHz            | 1.130     ||Jy                  |2.70E+09|  1.13E+00||Jy|1990PKS90.C...0000W|no uncertainty reported|    2700   MHz       | Broad-band measurement|04 11 58.2 +05 27 13 (B1950)| Integrated from scans|                                        |Homogenized from new and previously published data
35|2.5 GHz (ATCA)      | 1.20      || Jy                 |2.50E+09|  1.20E+00||Jy|2003PASJ...55..351T|no uncertainty reported|       2.5 GHz       | Broad-band measurement|| Flux integrated from map|                                        |From new raw data
36|1410 MHz            | 1.760     ||Jy                  |1.41E+09|  1.76E+00||Jy|1990PKS90.C...0000W|no uncertainty reported|    1410   MHz       | Broad-band measurement|04 11 58.2 +05 27 13 (B1950)| Integrated from scans|                                        |Homogenized from new and previously published data
37|1.4 GHz (ATCA)      | 1.86      || Jy                 |1.40E+09|  1.86E+00||Jy|2003PASJ...55..351T|no uncertainty reported|       1.4 GHz       | Broad-band measurement|| Flux integrated from map|                                        |From new raw data
38|1.40 GHz            | 2676      ||milliJy             |1.40E+09|  2.68E+00||Jy|1992ApJS...79..331W|no uncertainty reported|1.4        GHz       | Broad-band measurement|041158.7 +052718 (B1950)| Flux integrated from map|                                        |From new raw data
39|1.4GHz  (VLA)       | 2087.1    |+/-73.6 |milliJy             |1.40E+09|  2.09E+00|+/-7.36E-02|Jy|1998AJ....115.1693C|uncertainty|    1.40   GHz       | Broad-band measurement|04 14 37.75 +05 34 43.2 (J2000)| Flux integrated from map|High peak                               |From new raw data
40|635 MHz             | 3.700     ||Jy                  |6.35E+08|  3.70E+00||Jy|1990PKS90.C...0000W|no uncertainty reported|     635   MHz       | Broad-band measurement|04 11 58.2 +05 27 13 (B1950)| Integrated from scans|                                        |Homogenized from new and previously published data
41|408 MHz             | 3.09      |+/-0.15 |Jy                  |4.08E+08|  3.09E+00|+/-1.50E-01|Jy|1981MNRAS.194..693L|rms noise|408        MHz       | Broad-band measurement|041158.6 052707 (B1950)| Modelled datum|                                        |From new raw data; Corrected for contaminating sources
42|408 MHz             | 3.090     ||Jy                  |4.08E+08|  3.09E+00||Jy|1990PKS90.C...0000W|no uncertainty reported|     408   MHz       | Broad-band measurement|04 11 58.2 +05 27 13 (B1950)| Integrated from scans|                                        |Homogenized from new and previously published data
43|365 MHz (Texas)     | 2.916     |+/-0.036|Jy                  |3.65E+08|  2.92E+00|+/-3.60E-02|Jy|1996AJ....111.1945D|internal error|365        MHz       | Broad-band measurement; obtained by interpolation over frequency|041158.235 +052713.82 (B1950)| Integrated from scans|Model:P;MFlag:+;EFlag:+;LFlag:+.        |From new raw data
44|178 MHz             | 2.1       |+/-15.0%|Jy                  |1.78E+08|  2.10E+00|+/-3.15E-01|Jy|1967MmRAS..71...49G|uncertainty|178        MHz       | Broad-band measurement|041156.5 +052500 (B1950)| Integrated from scans|                                        |From new raw data; Uncorrected for known sources in beam
45|178 MHz             | 2.100     ||Jy                  |1.78E+08|  2.10E+00||Jy|1990PKS90.C...0000W|no uncertainty reported|     178   MHz       | Broad-band measurement|04 11 58.2 +05 27 13 (B1950)| Integrated from scans|                                        |Homogenized from new and previously published data
46|74 MHz (VLA)        | 0.88      |+/-0.14 | Jy                 |7.38E+07|  8.80E-01|+/-1.40E-01|Jy|2007AJ....134.1245C|rms uncertainty|    73.8   MHz       | Broad-band measurement|04 14 36.09 +05 34 39.4 (J2000)| Flux integrated from map|Corrected for clean bias                |From new raw data
