
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-04-04T09:22:48PDT



Photometric Data for SMM J221735.10+001533.3

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|I (Cousins)         | 23.58     |+/-0.08 |mag                 |3.79E+14|  9.43E-07|+/-7.21E-08|Jy|2004ApJ...616...71S|1 sigma|    7900   A         | Broad-band measurement| | Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
2|J (2MASS)           | 22.05     |+/-0.18 |mag                 |2.40E+14|  2.41E-06|+/-4.35E-07|Jy|2004ApJ...616...71S|1 sigma|    1.25   microns   | Broad-band measurement| | Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
3|K_s_ (2MASS)        | 20.28     |+/-0.14 |mag                 |1.38E+14|  5.15E-06|+/-7.09E-07|Jy|2004ApJ...616...71S|1 sigma|    2.17   microns   | Broad-band measurement| | Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
4|3.6 microns (IRAC)  | 4.3       |+/-0.5  |microJy             |8.44E+13|  4.30E-06|+/-5.00E-07|Jy|2009ApJ...699.1610H|uncertainty|     3.550 microns   | Broad-band measurement|22 17 35.16 +00 15 37.2 (J2000)| Flux in fixed aperture|                                        |From new raw data
5|4.5 microns (IRAC)  | 6.2       |+/-0.8  |microJy             |6.67E+13|  6.20E-06|+/-8.00E-07|Jy|2009ApJ...699.1610H|uncertainty|     4.493 microns   | Broad-band measurement|22 17 35.16 +00 15 37.2 (J2000)| Flux in fixed aperture|                                        |From new raw data
6|5.8 microns (IRAC)  | |<5.7       |microJy             |5.23E+13| |5.70E-06|Jy|2009ApJ...699.1610H|3 sigma|     5.731 microns   | Broad-band measurement|22 17 35.16 +00 15 37.2 (J2000)| Flux in fixed aperture|                                        |From new raw data
7|PAH 6.2 (Spitzer)   | |<0.77E-15  |erg/s/cm^2^         |4.84E+13| |1.59E-06|Jy|2009ApJ...699..667M|3rms uncertainty|       6.2 microns   | Line measurement; flux integrated over line; lines measured in emission|22 17 35.15 +00 15 37.2 (J2000)| Flux integrated from map|                                        |From new raw data
8|PAH 7.7 (Spitzer)   | |<0.37E-15  |erg/s/cm^2^         |3.89E+13|  7.25E-06|9.51E-07|Jy|2009ApJ...699..667M|3rms uncertainty|       7.7 microns   | Line measurement; flux integrated over line; lines measured in emission|22 17 35.15 +00 15 37.2 (J2000)| Flux integrated from map|                                        |From new raw data
9|8.0 microns (IRAC)  | 8.9       |+/-1.3  |microJy             |3.85E+13|  8.90E-06|+/-1.30E-06|Jy|2009ApJ...699.1610H|uncertainty|     7.782 microns   | Broad-band measurement|22 17 35.16 +00 15 37.2 (J2000)| Flux in fixed aperture|                                        |From new raw data
10|24 microns (MIPS)   | |<112.0     |microJy             |1.27E+13| |1.12E-04|Jy|2009ApJ...699.1610H|3 sigma|     23.68 microns   | Broad-band measurement|221735.15 +001537.2 (J2000)| Flux in fixed aperture|                                        |From new raw data
11|850 microns (SCUBA) | 6.3       |+/-1.3  |milliJy             |3.53E+11|  6.30E-03|+/-1.30E-03|Jy|2005ApJ...622..772C|uncertainty|     850   microns   | Broad-band measurement|221735.15 +001537.2 (J2000)| Flux integrated from map|                                        |From new raw data
12|CO(3-2) line (IRAM) | 0.8       |+/-0.2  |Jy km s^-1^         |3.46E+11|  1.59E-07|+/-3.97E-08|Jy|2005MNRAS.359.1165G|uncertainty|   3.099             | Line measurement; flux integrated over line; lines measured in emission|22 17 35.20 +00 15 37.6 (J2000)| Flux integrated from map|                                        |From new raw data
