
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-07-10T13:42:15PDT



Photometric Data for SPT-SJ214654-5507.8

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|3.6 microns (IRAC) |           |<0.0200|mJy             |8.44E+13||0.00200E-03|Jy|2011ApJ...728L...4H|3sigma uncertainty|     3.550 microns   | Broad-band measurement|09 13 05.0 -00 53 43 (J2000)| Flux in fixed aperture|                                        |From new raw data
2|4.5 microns (IRAC) |           |<0.0329|mJy             |6.67E+13||0.0329E-03|Jy|2011ApJ...728L...4H|3sigma uncertainty|     4.493 microns   | Broad-band measurement|09 13 05.0 -00 53 43 (J2000)| Flux in fixed aperture|                                        |From new raw data
3|100 microns (PACS) | 49.0      |+/-3.0  |mJy             |2.998e+12|49.0E-03|+/-3.0E-03             |Jy|2005MNRAS.358..149P|uncertainty|     850   microns   | Broad-band measurement|12 37 11.7 +62 22 12 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
4|160 microns (PACS) | 196.0    |+/-22.0 |mJy                |1.874e+12|196.0E-03|+/-25.0E-03  |Jy |2.40e+01          |3sigma|-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
5|250 microns (SPIRE)| 350.      |+/-25.0 |mJy             |1.199e+12| 350.0E-03|+/-25.0e-03 |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
5|250 microns (SPIRE)| 346.      |+/-36.0 |mJy             |1.199e+12| 346.0E-03|+/-36.0e-03 |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
6|350 microns (SPIRE)| 332.      |+/-23.  |mJy             |8.565e+11|332.E-03 |+/-23.0e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
6|350 microns (SPIRE)| 339.      |+/-35.  |mJy             |8.565e+11|339.E-03 |+/-35.0e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
1|350 microns (SABOCA) | 380.0 | 103. |milliJy      |8.56550e+11| 380.0E-3   |103.E-3 |Jy|2007MNRAS.376.1073Z|no uncertainty reported|     850   microns   | Broad-band measurement|02 39 51.9 -01 35 55 (J2000)| Flux integrated from map|S/N = 19.9                              |From reprocessed raw data
8|500 microns (SPIRE) | 269.     |+/-19. |mJy             |5.996e+11|269.0E-03 |+/-19.0e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
8|500 microns (SPIRE) | 257.     |+/-28. |mJy             |5.996e+11|257.0E-03 |+/-28.0e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
1|870 microns (LABOCA)| 101.0     |+/-7  |milliJy             |3.45E+11|  101.0E-03|+/-7.0E-03|Jy|2009ApJ...707.1201W|uncertainty|       870 microns   | Broad-band measurement|03 32 29.33 -27 56 19.3 (J2000)| Flux integrated from map|S/N = 4.6                               |From new raw data
1|870 microns (LABOCA)| 100.0     |+/-17  |milliJy             |3.45E+11|  100.0E-03|+/-17.0E-03|Jy|2009ApJ...707.1201W|uncertainty|       870 microns   | Broad-band measurement|03 32 29.33 -27 56 19.3 (J2000)| Flux integrated from map|S/N = 4.6                               |From new raw data
1|1.4 mm (SPT)        | 22.8     |+/-4.6 |milliJy             |2.20E+11|  22.8E-03|+/-4.6E-03|Jy|2010ApJ...719..763V|uncertainty|       1.4 mm        | Broad-band measurement|74.804 -59.708 (J2000)| Flux integrated from map|De-boosted flux; S/N = 7.05             |From new raw data
1|1.4 mm (SPT)        | 24.5     |+/-5.8 |milliJy             |2.20E+11|  24.5E-03|+/-5.8E-03|Jy|2010ApJ...719..763V|uncertainty|       1.4 mm        | Broad-band measurement|74.804 -59.708 (J2000)| Flux integrated from map|De-boosted flux; S/N = 7.05             |From new raw data
3|2.0 mm (SPT)        | 6.0     |+/-1.3 |milliJy             |1.50E+11|  6.0E-03|+/-1.3E-03|Jy|2010ApJ...719..763V|uncertainty|       2.0 mm        | Broad-band measurement|74.804 -59.708 (J2000)| Flux integrated from map|De-boosted flux; S/N = 6.20             |From new raw data
3|2.0 mm (SPT)        | 5.5     |+/-1.5 |milliJy             |1.50E+11|  5.5E-03|+/-1.5E-03|Jy|2010ApJ...719..763V|uncertainty|       2.0 mm        | Broad-band measurement|74.804 -59.708 (J2000)| Flux integrated from map|De-boosted flux; S/N = 6.20             |From new raw data
1|3.0mm (ALMA)        | 1.13 | 0.18 |milliJy            |1.0E+11| 1.13E-3 |0.18E-3 |Jy|2007MNRAS.376.1073Z|no uncertainty reported|     850   microns   | Broad-band measurement|02 39 51.9 -01 35 55 (J2000)| Flux integrated from map|S/N = 19.9                              |From reprocessed raw data
3|31.9GHz (ATCA)      | 140.0   |+/-20.0|microJy             |31.9E+09|140.0E-06|+/-20.0E-06|Jy|2010ApJ...719..763V|3sigma uncertainty|       2.0 mm        | Broad-band measurement|74.804 -59.708 (J2000)| Flux integrated from map|De-boosted flux; S/N = 6.20             |From new raw data
