
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-07-08T02:35:43PDT



Photometric Data for GOODS J123620.96+620714.6

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|B F435W (HST/ACS) AB      | 23.860    ||mag                 |6.98E+14|  1.04E-06||Jy|2007ApJ...660...81M|no uncertainty reported|    4297   A         | Broad-band measurement|12 36 20.943 +62 07 14.36 (J2000)| Flux integrated from map|                                        |From reprocessed raw data; Corrected for contaminatingsources
2|B (Subaru) AB       | 24.61     ||mag                 |6.77E+14|  5.20E-07||Jy|2006ApJ...653.1027W|no uncertainty reported| 4427.60   A         | Broad-band measurement|189.087262 62.120656 (J2000)| Flux in fixed aperture|3" diameter aperture                    |Averaged from previously published data
3|V (HST/ACS) AB      | 23.287    ||mag                 |5.08E+14|  1.76E-06||Jy|2007ApJ...660...81M|no uncertainty reported|    5907   A         | Broad-band measurement|12 36 20.943 +62 07 14.36 (J2000)| Flux integrated from map|                                        |From reprocessed raw data; Corrected for contaminatingsources
4|R (Keck II) AB      | 23.88     || mag                |4.62E+14|  1.02E-06||Jy|2004AJ....127.3121W|no uncertainty reported|   648.7   A         | Broad-band measurement|12 36 20.943 +62 07 14.36 (J2000)| Total flux|                                        |From new raw data
5|R (Subaru) AB       | 23.45     ||mag                 |4.59E+14|  1.51E-06||Jy|2006ApJ...653.1027W|no uncertainty reported| 6534.16   A         | Broad-band measurement|189.087262 62.120656 (J2000)| Flux in fixed aperture|3" diameter aperture                    |Averaged from previously published data
6|i F775W (HST/ACS) AB      | 22.504    ||mag                 |3.86E+14|  3.62E-06||Jy|2007ApJ...660...81M|no uncertainty reported|    7764   A         | Broad-band measurement|12 36 20.943 +62 07 14.36 (J2000)| Flux integrated from map|                                        |From reprocessed raw data; Corrected for contaminatingsources
7|I (Subaru) AB       | 22.81     ||mag                 |3.76E+14|  2.73E-06||Jy|2006ApJ...653.1027W|no uncertainty reported| 7975.89   A         | Broad-band measurement|189.087262 62.120656 (J2000)| Flux in fixed aperture|3" diameter aperture                    |Averaged from previously published data
8|z F850LP (HST/ACS) AB      | 21.764    ||mag                 |3.17E+14|  7.15E-06||Jy|2007ApJ...660...81M|no uncertainty reported|    9445   A         | Broad-band measurement|12 36 20.943 +62 07 14.36 (J2000)| Flux integrated from map|                                        |From reprocessed raw data; Corrected for contaminatingsources
9|HK' (QUIRC) AB      | 21.13     |+/-0.30 |mag                 |1.58E+14|  1.28E-05|+/-3.54E-06|Jy|2006ApJ...653.1027W|uncertainty|18947.38   A         | Broad-band measurement|189.087262 62.120656 (J2000)| Flux in fixed aperture|3" diameter aperture                    |Averaged from previously published data
10|24 microns (MIPS)   | 446.3     |+/-6.6  |microJy             |1.27E+13|  4.46E-04|+/-6.60E-06|Jy|2011A&A...528A..35M|uncertainty|     23.68 microns   | Broad-band measurement|12 36 20.94 +62 07 14.15 (J2000)| Flux integrated from map|                                        |From new raw data
1|24 microns (MIPS)   | 0.447     |+/-0.010 |mJy            |1.27E+13|0.447E-03|+/-0.010E-03|Jy|2009ApJ...694.1517D|1rms uncertainty|     23.68 microns   | Broad-band measurement|12 37 11.89 +62 22 11.8 (J2000)| Flux integrated from map|                                        |From new raw data
11|70 microns (MIPS)   | 5.8       |+/-0.3  |milliJy             |4.20E+12|  5.80E-03|+/-3.00E-04|Jy|2011A&A...528A..35M|uncertainty|     71.42 microns   | Broad-band measurement|12 36 20.94 +62 07 14.15 (J2000)| Flux integrated from map|                                        |From new raw data
2|70 microns (MIPS)   | 5.3       |+/-0.7   |mJy            |4.20E+12|5.3E-03  |+/-0.7E-03|Jy|2009ApJ...699.1610H|3 sigma|     71.42 microns   | Broad-band measurement|221804.42 +002154.4 (J2000)| Flux in fixed aperture|                                        |From new raw data
12|1.4 GHz (VLA)             | 90.4      |+/-9.6  |microJy             |1.40E+09|  9.04E-05|+/-9.60E-06|Jy|2000ApJ...533..611R|1 sigma|1.4        GHz       | Broad-band measurement; broad-band flux derived by integration over spectrum; synthetic band|123620.983 +620713.87 (J2000)| Flux integrated from map; Pointing and beam filling|                                        |From new raw data; Corrected for contaminating sources
