
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-05-27T06:38:15PDT



Photometric Data for SHADES J021725-045937

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|B (SUBARU) AB        | 24.38    |+/-0.032|mag   |6.69E+14|  6.43E-07|+/-1.89E-08|Jy|2008MNRAS.387..247C|uncertainty|      4478 A         | Broad-band measurement|34.354730 -4.992860 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
2|V (SUBARU) AB        | 24.30    |+/-0.029|mag   |5.46E+14|  6.92E-07|+/-1.85E-08|Jy|2008MNRAS.387..247C|uncertainty|      5493 A         | Broad-band measurement|34.354730 -4.992860 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
3|R (SUBARU) AB        | 24.09    |+/-0.030|mag   |4.58E+14|  8.40E-07|+/-2.32E-08|Jy|2008MNRAS.387..247C|uncertainty|      6550 A         | Broad-band measurement|34.354730 -4.992860 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
4|i' (SUBARU) AB       | 23.97    |+/-0.032|mag   |3.89E+14|  9.38E-07|+/-2.76E-08|Jy|2008MNRAS.387..247C|uncertainty|      7709 A         | Broad-band measurement|34.354730 -4.992860 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
5|z' (SUBARU) AB       | 23.66    |+/-0.029|mag   |3.31E+14|  1.25E-06|+/-3.33E-08|Jy|2008MNRAS.387..247C|uncertainty|      9054 A         | Broad-band measurement|34.354730 -4.992860 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
7|3.6 microns (IRAC)  | 2.5993E+01|+/-1.0118E+00|microJy             |8.44E+13|  2.60E-05|+/-1.01E-06|Jy|2013SSTSLC4.2....0C|uncertainty|3.55       microns   | Broad-band measurement|| Flux in fixed aperture|5.8" aperture                           |From new raw data
8|3.6 microns (IRAC)  | 3.2925E+01|+/-1.8243E-01|microJy             |8.44E+13|  3.29E-05|+/-1.82E-07|Jy|2013SSTSLC4.2....0C|uncertainty|3.55       microns   | Broad-band measurement|| Flux in fixed aperture|5.8" aperture                           |From new raw data
12|4.5 microns (IRAC)  | 2.6923E+01|+/-1.6337E+00|microJy             |6.67E+13|  2.69E-05|+/-1.63E-06|Jy|2013SSTSLC4.2....0C|uncertainty|4.493      microns   | Broad-band measurement|| Flux in fixed aperture|5.8" aperture                           |From new raw data
13|4.5 microns (IRAC)  | 3.6368E+01|+/-2.2095E-01|microJy             |6.67E+13|  3.64E-05|+/-2.21E-07|Jy|2013SSTSLC4.2....0C|uncertainty|4.493      microns   | Broad-band measurement|| Flux in fixed aperture|5.8" aperture                           |From new raw data
6|4.5 microns (IRAC)   | 21.35    |+/-1.08 |uJy   |6.67E+13|  2.14E-05|+/-1.08E-06|Jy|2008MNRAS.387..247C|uncertainty|     4.493 microns   | Broad-band measurement|34.354730 -4.992860 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
16|5.8 microns (IRAC)  | 3.2512E+01|+/-8.2667E-01|microJy             |5.23E+13|  3.25E-05|+/-8.27E-07|Jy|2013SSTSLC4.2....0C|uncertainty|5.731      microns   | Broad-band measurement|| Flux in fixed aperture|5.8" aperture                           |From new raw data
18|5.8 microns (IRAC)  | 6.1606E+01|+/-6.6572E+00|microJy             |5.23E+13|  6.16E-05|+/-6.66E-06|Jy|2013SSTSLC4.2....0C|uncertainty|5.731      microns   | Broad-band measurement|| Flux in fixed aperture|5.8" aperture                           |From new raw data
21|8.0 microns (IRAC)  | 3.2766E+01|+/-1.1327E+00|microJy             |3.81E+13|  3.28E-05|+/-1.13E-06|Jy|2013SSTSLC4.2....0C|uncertainty|7.872      microns   | Broad-band measurement|| Flux in fixed aperture|5.8" aperture                           |From new raw data
7|15 microns (AKARI)   | 105      |+/-20   |uJy   |1.92E+13|  1.05E-04|+/-2.00E-05|Jy|2010A&A...514A..10S|uncertainty|     15.58 microns   | Broad-band measurement| | Flux in fixed aperture|                                        |From new raw data
8|24 microns (Spitzer/MIPS) | 195.0    |+/-47.0 |uJy   |1.27E+13|  1.95E-04|+/-4.70E-05|Jy|2007MNRAS.380..199I|rms uncertainty|     23.68 microns   | Broad-band measurement|02 17 25.16 -04 59 35.0 (J2000)| Flux integrated from map|                                        |Averaged from previously published data
9|24 microns (MIPS)    | 212.34   |+/-15.22|uJy   |1.27E+13|  2.12E-04|+/-1.52E-05|Jy|2008MNRAS.387..247C|uncertainty|     23.68 microns   | Broad-band measurement|34.354730 -4.992860 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
25|24 microns (MIPS)   | 2.2110E+02|+/-1.0142E+01|microJy             |1.27E+13|  2.21E-04|+/-1.01E-05|Jy|2013SSTSLC4.2....0C|uncertainty|23.68      microns   | Broad-band measurement|| Modelled datum|PSF fit                                 |From new raw data
26|24 microns (MIPS)   | 1.7652E+02|+/-5.1917E+01|microJy             |1.27E+13|  1.77E-04|+/-5.19E-05|Jy|2013SSTSLC4.2....0C|uncertainty|23.68      microns   | Broad-band measurement|| Modelled datum|PSF fit                                 |From new raw data
27|24 microns (MIPS)   | 2.3731E+02|+/-9.4247E+00|microJy             |1.27E+13|  2.37E-04|+/-9.42E-06|Jy|2013SSTSLC4.2....0C|uncertainty|23.68      microns   | Broad-band measurement|| Flux in fixed aperture|14.7" aperture                          |From new raw data
28|24 microns (MIPS)   | 1.9630E+02|+/-4.7772E+01|microJy             |1.27E+13|  1.96E-04|+/-4.78E-05|Jy|2013SSTSLC4.2....0C|uncertainty|23.68      microns   | Broad-band measurement|| Flux in fixed aperture|14.7" aperture                          |From new raw data
10|250 microns (SPIRE) | 21.7     |+/-3.6  |mJy   |1.199e+12| 21.7E-03|+/-3.6E-03  |Jy|Reference          |uncertainty       | | | | |
11|350 microns (SPIRE) | 22.2     |+/-4.2  |mJy   |8.57e+11|  22.2E-03|+/-4.2E-03  |Jy|Reference          |uncertainty       | | | | |
12|350 microns (CSO/SHARC-II)   | 31.1     |+/-15.0 |mJy   |8.57E+11|  3.11E-02|+/-1.50E-02|Jy|2008MNRAS.384.1597C|uncertainty|       350 microns   | Broad-band measurement| | Flux integrated from map|Corrected for flux boosting             |From new raw data
13|500 microns (SPIRE) | 17.0     |+/-4.8  |mJy   |5.996e+11| 17.0E-03|+/-4.8E-03  |Jy|Reference          |uncertainty       | | | | |
14|850 microns (SCUBA) | 4.5      |+/-2.2  |mJy   |3.53E+11|  4.50E-03|+/-2.20E-03|Jy|2007MNRAS.380..199I|rms uncertainty|       850 microns   | Broad-band measurement|02 17 25.117 -04 59 37.44 (J2000)| Flux integrated from map|                                        |Averaged from previously published data
15|850 microns (SCUBA) | 4.5      |+/-1.9  |mJy   |3.53E+11|  4.50E-03|+/-1.90E-03|Jy|2008MNRAS.387..247C|uncertainty|       850 microns   | Broad-band measurement|34.354730 -4.992860 (J2000)| Flux integrated from map|                                        |Averaged from previously published data
16|1.4 GHz (VLA)       | 56.8     |+/-10.0 |uJy   |1.40E+09|  5.68E-05|+/-1.00E-05|Jy|2007MNRAS.380..199I|rms uncertainty|       1.4 GHz       | Broad-band measurement|02 17 25.101 -04 59 33.77 (J2000)| Flux integrated from map|                                        |From new raw data
