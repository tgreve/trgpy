
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-06-17T13:44:57PDT



Photometric Data for GOODS J123711.48+622155.8

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|U (KPNO) AB         ||>26.7      |mag                 |8.44E+14||7.59E-08|Jy|2009A&A...500..705M|3 sigma|      3552 A         | Broad-band measurement|12 37 11.5 +62 21 55.8 (J2000)| Flux in fixed aperture|                                        |From new raw data
2|B (HST) AB          ||>26.3      |mag                 |6.98E+14||1.10E-07|Jy|2009A&A...500..705M|3 sigma|      4297 A         | Broad-band measurement|12 37 11.5 +62 21 55.8 (J2000)| Flux in fixed aperture|                                        |From new raw data
3|F435W (HST) AB      | 28.90     |+/-1.70 |mag                 |6.98E+14|  1.00E-08|+/-1.57E-08|Jy|2011ApJ...738...69S|uncertainty|      4297 A         | Broad-band measurement|12 37 11.48 +62 21 55.83 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
4|V (HST) AB          | 25.010    ||mag                 |5.08E+14|  3.60E-07||Jy|2009A&A...500..705M|no uncertainty reported|      5907 A         | Broad-band measurement|12 37 11.5 +62 21 55.8 (J2000)| Flux in fixed aperture|                                        |From new raw data
5|F606W (HST) AB      | 25.04     |+/-0.07 |mag                 |5.08E+14|  3.50E-07|+/-2.26E-08|Jy|2011ApJ...738...69S|uncertainty|      5907 A         | Broad-band measurement|12 37 11.48 +62 21 55.83 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
6|R (Keck II) AB      | 24.55     || mag                |4.62E+14|  5.50E-07||Jy|2004AJ....127.3121W|no uncertainty reported|   648.7   A         | Broad-band measurement|12 37 11.477 +62 21 55.35 (J2000)| Total flux|                                        |From new raw data
7|i (HST) AB          | 23.929    ||mag                 |3.86E+14|  9.74E-07||Jy|2009A&A...500..705M|no uncertainty reported|      7764 A         | Broad-band measurement|12 37 11.5 +62 21 55.8 (J2000)| Flux in fixed aperture|                                        |From new raw data
8|F775W (HST) AB      | 23.99     |+/-0.06 |mag                 |3.86E+14|  9.21E-07|+/-5.09E-08|Jy|2011ApJ...738...69S|uncertainty|      7764 A         | Broad-band measurement|12 37 11.48 +62 21 55.83 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
9|z (HST) AB          | 23.658    ||mag                 |3.17E+14|  1.25E-06||Jy|2009A&A...500..705M|no uncertainty reported|      9445 A         | Broad-band measurement|12 37 11.5 +62 21 55.8 (J2000)| Flux in fixed aperture|                                        |From new raw data
10|F850LP (HST) AB     | 23.66     |+/-0.05 |mag                 |3.17E+14|  1.25E-06|+/-5.75E-08|Jy|2011ApJ...738...69S|uncertainty|      9445 A         | Broad-band measurement|12 37 11.48 +62 21 55.83 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
11|J (KPNO) AB         | 23.133    ||mag                 |2.40E+14|  2.03E-06||Jy|2009A&A...500..705M|no uncertainty reported|  1247.975 nm        | Broad-band measurement|12 37 11.5 +62 21 55.8 (J2000)| Flux in fixed aperture|                                        |From new raw data
12|J (CFHT) AB         | 23.61     |+/-0.09 |mag                 |2.40E+14|  1.31E-06|+/-1.08E-07|Jy|2011ApJ...738...69S|uncertainty|      1.25 microns   | Broad-band measurement|12 37 11.48 +62 21 55.83 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
13|H (KPNO) AB         | 23.167    ||mag                 |1.83E+14|  1.96E-06||Jy|2009A&A...500..705M|no uncertainty reported|    1635.6 nm        | Broad-band measurement|12 37 11.5 +62 21 55.8 (J2000)| Flux in fixed aperture|                                        |From new raw data
14|K_s(KPNO) AB        | 23.125    ||mag                 |1.40E+14|  2.04E-06||Jy|2009A&A...500..705M|no uncertainty reported|    2147.5 nm        | Broad-band measurement|12 37 11.5 +62 21 55.8 (J2000)| Flux in fixed aperture|                                        |From new raw data
15|K (CFHT) AB         | 22.92     |+/-0.10 |mag                 |1.39E+14|  2.47E-06|+/-2.27E-07|Jy|2011ApJ...738...69S|uncertainty|      2.15 microns   | Broad-band measurement|12 37 11.48 +62 21 55.83 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
16|3.6 microns IRAC AB | 22.352    ||mag                 |8.44E+13|  4.16E-06||Jy|2009A&A...500..705M|no uncertainty reported|     3.550 microns   | Broad-band measurement|12 37 11.5 +62 21 55.8 (J2000)| Flux in fixed aperture|                                        |From new raw data
17|3.6 microns IRAC AB | 22.34     |+/-0.06 |mag                 |8.44E+13|  4.21E-06|+/-2.33E-07|Jy|2011ApJ...738...69S|uncertainty|     3.550 microns   | Broad-band measurement|12 37 11.48 +62 21 55.83 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
18|4.5 microns IRAC AB | 22.714    ||mag                 |6.67E+13|  2.98E-06||Jy|2009A&A...500..705M|no uncertainty reported|     4.493 microns   | Broad-band measurement|12 37 11.5 +62 21 55.8 (J2000)| Flux in fixed aperture|                                        |From new raw data
19|4.5 microns IRAC AB | 22.73     |+/-0.06 |mag                 |6.67E+13|  2.94E-06|+/-1.62E-07|Jy|2011ApJ...738...69S|uncertainty|     4.493 microns   | Broad-band measurement|12 37 11.48 +62 21 55.83 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
20|5.8 microns IRAC AB | 22.64     |+/-0.17 |mag                 |5.23E+13|  3.19E-06|+/-5.00E-07|Jy|2011ApJ...738...69S|uncertainty|     5.731 microns   | Broad-band measurement|12 37 11.48 +62 21 55.83 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
21|8.0 microns IRAC AB | 22.414    ||mag                 |3.81E+13|  3.93E-06||Jy|2009A&A...500..705M|no uncertainty reported|     7.872 microns   | Broad-band measurement|12 37 11.5 +62 21 55.8 (J2000)| Flux in fixed aperture|                                        |From new raw data
22|8.0 microns IRAC AB | 22.33     |+/-0.13 |mag                 |3.81E+13|  4.25E-06|+/-5.08E-07|Jy|2011ApJ...738...69S|uncertainty|     7.872 microns   | Broad-band measurement|12 37 11.48 +62 21 55.83 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
23|24 microns (MIPS)   | 52.6      |+/-2.2  |microJy             |1.27E+13|  5.26E-05|+/-2.20E-06|Jy|2011A&A...528A..35M|uncertainty|     23.68 microns   | Broad-band measurement|12 37 11.49 +62 21 55.50 (J2000)| Flux integrated from map|                                        |From new raw data
24|24 microns MIPS AB  | 19.934    ||mag                 |1.27E+13|  3.86E-05||Jy|2009A&A...500..705M|no uncertainty reported|     23.68 microns   | Broad-band measurement|12 37 11.5 +62 21 55.8 (J2000)| Flux in fixed aperture|                                        |From new raw data
25|70 microns (MIPS)   ||<4.7       |milliJy             |4.20E+12||4.70E-03|Jy|2011A&A...528A..35M|no uncertainty reported|     71.42 microns   | Broad-band measurement|12 37 11.49 +62 21 55.50 (J2000)| Flux integrated from map|                                        |From new raw data
