
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-07-10T13:42:15PDT



Photometric Data for SPT-SJ214654-5507.8

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|3.6 microns (IRAC) | 0.0020   |+/-0.0006|mJy             |8.44E+13|0.0020E-03|+/-0.0006E-03|Jy|2011ApJ...728L...4H|3sigma uncertainty|     3.550 microns   | Broad-band measurement|09 13 05.0 -00 53 43 (J2000)| Flux in fixed aperture|                                        |From new raw data
2|4.5 microns (IRAC) | 0.0035   |+/-0.0004|mJy             |6.67E+13|0.0035E-03|+/-0.0004E-03|Jy|2011ApJ...728L...4H|3sigma uncertainty|     4.493 microns   | Broad-band measurement|09 13 05.0 -00 53 43 (J2000)| Flux in fixed aperture|                                        |From new raw data
3|100 microns (PACS) | 9.0      |+/-2.0  |mJy             |2.998e+12|9.0E-03|+/-2.0E-03             |Jy|2005MNRAS.358..149P|uncertainty|     850   microns   | Broad-band measurement|12 37 11.7 +62 22 12 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
4|160 microns (PACS) |          |<28.0 |mJy                |1.874e+12|         |28.0E-03  |Jy |2.40e+01          |3sigma|-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
5|250 microns (SPIRE)| 72.      |+/-9.0 |mJy             |1.199e+12| 72.0E-03|+/-9.0e-03 |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
6|350 microns (SPIRE)| 115.      |+/-10.  |mJy             |8.565e+11|115.E-03 |+/-10.0e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
8|500 microns (SPIRE) | 121.     |+/-11. |mJy             |5.996e+11|121.0E-03 |+/-11.0e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
1|870 microns (LABOCA)| 61.0     |+/-5  |milliJy             |3.45E+11|  61.0E-03|+/-5.0E-03|Jy|2009ApJ...707.1201W|uncertainty|       870 microns   | Broad-band measurement|03 32 29.33 -27 56 19.3 (J2000)| Flux integrated from map|S/N = 4.6                               |From new raw data
1|1.4 mm (SPT)        | 20.3     |+/-4.6 |milliJy             |2.20E+11|  20.3E-03|+/-4.6E-03|Jy|2010ApJ...719..763V|uncertainty|       1.4 mm        | Broad-band measurement|74.804 -59.708 (J2000)| Flux integrated from map|De-boosted flux; S/N = 7.05             |From new raw data
3|2.0 mm (SPT)        | 5.8     |+/-1.3 |milliJy             |1.50E+11|  5.8E-03|+/-1.3E-03|Jy|2010ApJ...719..763V|uncertainty|       2.0 mm        | Broad-band measurement|74.804 -59.708 (J2000)| Flux integrated from map|De-boosted flux; S/N = 6.20             |From new raw data
3|47.5GHz (ATCA)      | 140.0   |+/-40.0|microJy             |47.5E+09|140.0E-06|+/-40.0E-06|Jy|2010ApJ...719..763V|3sigma uncertainty|       2.0 mm        | Broad-band measurement|74.804 -59.708 (J2000)| Flux integrated from map|De-boosted flux; S/N = 6.20             |From new raw data
