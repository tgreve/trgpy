

Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.


queryDateTime:2009-11-03T15:07:35PST








No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|U (WHT)            |       |>27.2  |mag                 |8.48549e+14|  |4.78628e-08|Jy|2004ApJ...616...71S|3sigma uncertainty|    1.25   microns   | Broad-band measurement| | Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
1|g (WHT)            |       |>27.3  |mag                 |6.17874e+14|  |4.78628e-08 |Jy|2004ApJ...616...71S|3sigma uncertainty|    1.25   microns   | Broad-band measurement| | Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
1|R (Cousins) AB      | 27.0      |+/-0.3  |mag                 |4.72E+14|  5.755e-08|+/-1.15549e-08 |Jy|2004ApJ...616...71S|sigma uncertainty|    1.25   microns   | Broad-band measurement| | Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
2|HST/ACS F814W AB    | 26.0      |+/-0.2  |mag                 |3.78E+14|  1.446e-07   |+/-2.924e-08|Jy|2004A&A...421..847Z|no uncertainty reported|    7924   A         | Broad-band measurement| | Flux in fixed aperture|3" aperture                             |From reprocessed raw data
3|J (Bessel) AB       | 23.92     |+/-0.2  |mag                 |2.40E+14|  9.818e-07|+/-1.986e-07|Jy|2004ApJ...616...71S|sigma uncertainty|    1.25   microns   | Broad-band measurement| | Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
4|K (Bessel) AB       | 22.3      |+/-0.2  |mag                 |1.38E+14|  4.365e-06|+/-8.830e-07|Jy|2004ApJ...616...71S|sigma uncertainty|    1.25   microns   | Broad-band measurement| | Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
5|IRAC 4.5um          | 21.9      |+/-0.2  |microJy            |6.67E+13|  6.310e-06|+/-1.831e-08|Jy|1996AJ....111.1431B|uncertainty|1.49       GHz       | Broad-band measurement| | Peak flux|                                        |From new raw data
6|MIPS 24um           | 160.1     |+/-5.0  |microJy             |1.27E+13|  160.1E-06  |+/-5.0E-06 |Jy|1996AJ....111.1431B|uncertainty|1.49       GHz       | Broad-band measurement| | Peak flux|                                        |From new raw data
7|SMA 870um           |           |<3.3    |milliJy             |340.0E+09|            |3.3E-03 |Jy|1996AJ....111.1431B|3sigma uncertainty|1.49       GHz       | Broad-band measurement| | Peak flux|                                        |From new raw data
