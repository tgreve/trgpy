
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-07-10T08:38:10PDT



Photometric Data for LESS 073

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|2-10 keV (Chandra)  | 7.24E-16  ||erg cm^-2^ s^-1^    |1.45E+18|  4.99E-11||Jy|2006A&A...451..457T|no uncertainty reported|       6   keV       | Broad-band measurement|| Flux integrated from map|                                        |From reprocessed raw data; NED frequency assigned tomid-point of band in keV
2|2-10 keV (Chandra)  | 6.8E-16   |+/-2.4E-16|erg/cm^2^/s         |1.45E+18|  4.69E-11|+/-1.66E-11|Jy|2011ApJ...730L..28G|uncertainty|     6.00  keV       | Broad-band measurement|03 32 29.29 -27 56 19.5 (J2000)| Flux in fixed aperture|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
3|2-8 keV (Chandra)   ||<7.6E-16   |erg s^-1^ cm^-2^    |1.21E+18||6.28E-11|Jy|2007A&A...461...39F|3sigma no uncertainty reported|       5   keV       | Broad-band measurement|03 32 29.29 -27 56 19.4 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data; NED frequencyassigned to mid-point of band in keV
4|2-8 keV (Chandra)   | 5.0E-16   ||erg/cm^2^/s         |1.21E+18|  4.13E-11||Jy|2011ApJS..195...10X|no uncertainty reported|      5.00 keV       | Broad-band measurement|03 32 29.27 -27 56 19.8 (J2000)| Modelled datum|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
5|0.5-8 keV (Chandra) | 5.0E-16   ||erg/cm^2^/s         |1.03E+18|  4.85E-11||Jy|2011ApJS..195...10X|no uncertainty reported|      4.25 keV       | Broad-band measurement|03 32 29.27 -27 56 19.8 (J2000)| Modelled datum|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
6|0.5-2 keV (Chandra) | 0.50E-16  ||erg s^-1^ cm^-2^    |3.02E+17|  1.66E-11||Jy|2007A&A...461...39F|no uncertainty reported|    1.25   keV       | Broad-band measurement|03 32 29.29 -27 56 19.4 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data; NED frequencyassigned to mid-point of band in keV
7|0.5-2 keV (Chandra) | 1.11E-16  ||erg cm^-2^ s^-1^    |3.02E+17|  3.68E-11||Jy|2006A&A...451..457T|no uncertainty reported|    1.25   keV       | Broad-band measurement|| Flux integrated from map|                                        |From reprocessed raw data; NED frequency assigned tomid-point of band in keV
8|0.5-2 keV (Chandra) | 4.2E-17   |+/-1.5E-17|erg/cm^2^/s         |3.02E+17|  1.39E-11|+/-4.97E-12|Jy|2011ApJ...730L..28G|uncertainty|     1.25  keV       | Broad-band measurement|03 32 29.29 -27 56 19.5 (J2000)| Flux in fixed aperture|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
9|0.5-2 keV (Chandra) ||<7.3E-17   |erg/cm^2^/s         |3.02E+17||2.42E-11|Jy|2011ApJS..195...10X|3sigma no uncertainty reported|      1.25 keV       | Broad-band measurement|03 32 29.27 -27 56 19.8 (J2000)| Modelled datum|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
10|0.5-2 keV (Chandra) | 1.0E-16   ||erg/cm^2^/s         |3.02E+17|  3.31E-11||Jy|2012A&A...537A..16F|no uncertainty reported|      1.25 keV       | Broad-band measurement|53.122036 -27.938740 (J2000)| Modelled datum|                                        |From reprocessed raw data; NED frequency assigned tomid-point of band in keV
11|U                   | 4.528E-03 |+/-1.908E-03|photons/m^2^/s/nm   |8.21E+14|  1.10E-07|+/-4.61E-08|Jy|2004A&A...421..913W|1 sigma| 365       nm        | Broad-band measurement|033229.289 -275619.36 (J2000)| Flux in fixed aperture|          0          01.5" aperture     |From new raw data
12|418 nm              | 3.663E-03 |+/-3.279E-03|photons/m^2^/s/nm   |7.17E+14|  1.02E-07|+/-9.08E-08|Jy|2004A&A...421..913W|1 sigma| 418       nm        | Broad-band measurement|033229.289 -275619.36 (J2000)| Flux in fixed aperture|          0          01.5" aperture     |From new raw data
13|F435W (HST/ACS) AB  ||>29.82     |mag                 |6.98E+14||4.29E-09|Jy|2004ApJ...600L.119C|3sigma no uncertainty reported|    4297   A         | Broad-band measurement|03 32 29.29 -27 56 19.3 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data; derived from a fluxin a different band and a color
14|F435W (HST) AB      ||>28.86     |mag                 |6.98E+14||1.04E-08|Jy|2010A&A...510A.109R|3sigma no uncertainty reported|      4297 A         | Broad-band measurement|03 32 29.29 -27 56 19.5 (J2000)| Flux in fixed aperture|Corrected to 6" circular aperture       |From reprocessed raw data
15|F435W (HST/ACS) AB  ||>29.84     |mag                 |6.98E+14||4.19E-09|Jy|2007A&A...461...39F|3sigma no uncertainty reported|    4297   A         | Broad-band measurement|03 32 29.29 -27 56 19.4 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data; derived from a fluxin a different band and a color
16|F435W (HST) AB      ||>28.90     |mag                 |6.98E+14||1.00E-08|Jy|2011ApJ...738...69S|3 sigma|      4297 A         | Broad-band measurement|03 32 29.29 -27 56 19.46 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
18|462 nm              | 2.213E-03 |+/-3.065E-03|photons/m^2^/s/nm   |6.49E+14|  6.78E-08|+/-9.38E-08|Jy|2004A&A...421..913W|1 sigma| 462       nm        | Broad-band measurement|033229.289 -275619.36 (J2000)| Flux in fixed aperture|          0          01.5" aperture     |From new raw data
19|486 nm              | 7.523E-04 |+/-3.904E-03|photons/m^2^/s/nm   |6.17E+14|  2.42E-08|+/-1.26E-07|Jy|2004A&A...421..913W|1 sigma| 486       nm        | Broad-band measurement|033229.289 -275619.36 (J2000)| Flux in fixed aperture|          0          01.5" aperture     |From new raw data
20|519 nm              | 5.132E-03 |+/-4.871E-03|photons/m^2^/s/nm   |5.78E+14|  1.76E-07|+/-1.68E-07|Jy|2004A&A...421..913W|1 sigma| 519       nm        | Broad-band measurement|033229.289 -275619.36 (J2000)| Flux in fixed aperture|          0          01.5" aperture     |From new raw data
21|V                   | 1.026E-03 |+/-1.651E-03|photons/m^2^/s/nm   |5.57E+14|  3.66E-08|+/-5.89E-08|Jy|2004A&A...421..913W|1 sigma| 538       nm        | Broad-band measurement|033229.289 -275619.36 (J2000)| Flux in fixed aperture|          0          01.5" aperture     |From new raw data
22|V                   | 27.545    |+/-1.000|mag                 |5.45E+14|  3.49E-08|+/-5.28E-08|Jy|2001A&A...377..442W|mean error|5500       A         | Broad-band measurement|033229.289 -275619.36 (J2000)| Corrected to total flux from single aperture measurement|                                        |From new raw data
23|572 nm              | 9.441E-04 |+/-3.514E-03|photons/m^2^/s/nm   |5.24E+14|  3.58E-08|+/-1.33E-07|Jy|2004A&A...421..913W|1 sigma| 572       nm        | Broad-band measurement|033229.289 -275619.36 (J2000)| Flux in fixed aperture|          0          01.5" aperture     |From new raw data
24|F606W (HST/ACS) AB  | 26.76     |+/-0.09 |mag                 |5.08E+14|  7.18E-08|+/-5.95E-09|Jy|2007ApJ...659...84S|uncertainty|    5907   A         | Broad-band measurement|03 32 29.29 -27 56 19.46 (J2000)| Corrected to total flux from single aperture measurement|                                        |From reprocessed raw data; Extinction-corrected for Milky Way
25|F606W (HST) AB      | 26.93     |+/-0.14 |mag                 |5.08E+14|  6.14E-08|+/-7.92E-09|Jy|2010A&A...510A.109R|uncertainty|      5907 A         | Broad-band measurement|03 32 29.29 -27 56 19.5 (J2000)| Flux in fixed aperture|Corrected to 6" circular aperture       |From reprocessed raw data
26|F606W (HST/ACS) AB  | 26.84     ||mag                 |5.08E+14|  6.64E-08||Jy|2007A&A...461...39F|no uncertainty reported|    5907   A         | Broad-band measurement|03 32 29.29 -27 56 19.4 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data; derived from a fluxin a different band and a color
27|F606W (HST/ACS) AB  | 26.82     ||mag                 |5.08E+14|  6.79E-08||Jy|2004ApJ...600L.119C|no uncertainty reported|    5907   A         | Broad-band measurement|03 32 29.29 -27 56 19.3 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data; derived from a fluxin a different band and a color
28|F606W (HST) AB      | 26.83     |+/-0.10 |mag                 |5.08E+14|  6.73E-08|+/-6.20E-09|Jy|2011ApJ...738...69S|uncertainty|      5907 A         | Broad-band measurement|03 32 29.29 -27 56 19.46 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
29|605 nm              | 2.178E-03 |+/-3.599E-03|photons/m^2^/s/nm   |4.96E+14|  8.73E-08|+/-1.44E-07|Jy|2004A&A...421..913W|1 sigma| 605       nm        | Broad-band measurement|033229.289 -275619.36 (J2000)| Flux in fixed aperture|          0          01.5" aperture     |From new raw data
30|R                   | 25.302    |+/-0.126|mag                 |4.68E+14|  2.33E-07|+/-2.87E-08|Jy|2001A&A...377..442W|mean error|6400       A         | Broad-band measurement|033229.289 -275619.36 (J2000)| Corrected to total flux from single aperture measurement|                                        |From new raw data
31|645 nm              | 1.796E-02 |+/-6.752E-03|photons/m^2^/s/nm   |4.65E+14|  7.68E-07|+/-2.89E-07|Jy|2004A&A...421..913W|1 sigma| 645       nm        | Broad-band measurement|033229.289 -275619.36 (J2000)| Flux in fixed aperture|          0          01.5" aperture     |From new raw data
32|R (total)           | 25.606    |+/-0.249|mag                 |4.63E+14|  2.08E-07|+/-4.77E-08|Jy|2004A&A...421..913W|1 sigma| 648       nm        | Broad-band measurement|033229.289 -275619.36 (J2000)| Flux integrated from map|          0          01.5" aperture     |From new raw data
33|R                   | 6.059E-03 |+/-4.764E-04|photons/m^2^/s/nm   |4.63E+14|  2.60E-07|+/-2.05E-08|Jy|2004A&A...421..913W|1 sigma| 648       nm        | Broad-band measurement|033229.289 -275619.36 (J2000)| Flux in fixed aperture|          0          01.5" aperture     |From new raw data
34|696 nm              | 1.715E-02 |+/-2.943E-03|photons/m^2^/s/nm   |4.31E+14|  7.91E-07|+/-1.36E-07|Jy|2004A&A...421..913W|1 sigma| 696       nm        | Broad-band measurement|033229.289 -275619.36 (J2000)| Flux in fixed aperture|          0          01.5" aperture     |From new raw data
35|753 nm              | 2.113E-02 |+/-4.959E-03|photons/m^2^/s/nm   |3.98E+14|  1.05E-06|+/-2.47E-07|Jy|2004A&A...421..913W|1 sigma| 753       nm        | Broad-band measurement|033229.289 -275619.36 (J2000)| Flux in fixed aperture|          0          01.5" aperture     |From new raw data
36|F775W (HST) AB      | 25.2020   || mag                |3.86E+14|  3.02E-07||Jy|2008A&A...478...83V|no uncertainty reported|      7764 A         | Broad-band measurement|033229.29 -275619.5 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data; derived from aflux in a different band and a color
37|F775W (HST) AB      | 25.12     |+/-0.04 |mag                 |3.86E+14|  3.25E-07|+/-1.20E-08|Jy|2010A&A...510A.109R|uncertainty|      7764 A         | Broad-band measurement|03 32 29.29 -27 56 19.5 (J2000)| Flux in fixed aperture|Corrected to 6" circular aperture       |From reprocessed raw data
38|F775W (HST/ACS) AB  | 25.17     ||mag                 |3.86E+14|  3.11E-07||Jy|2004ApJ...600L.119C|no uncertainty reported|    7764   A         | Broad-band measurement|03 32 29.29 -27 56 19.3 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data; derived from a fluxin a different band and a color
39|F775W (HST/ACS) AB  | 25.12     ||mag                 |3.86E+14|  3.25E-07||Jy|2006A&A...454..423V|no uncertainty reported|    7764   A         | Broad-band measurement|033229.29 -275619.5 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data; derived from aflux in a different band and a color
40|F775W (HST/ACS) AB  | 25.04     |+/-0.04 |mag                 |3.86E+14|  3.50E-07|+/-1.29E-08|Jy|2007ApJ...659...84S|uncertainty|    7764   A         | Broad-band measurement|03 32 29.29 -27 56 19.46 (J2000)| Corrected to total flux from single aperture measurement|                                        |From reprocessed raw data; Extinction-corrected for Milky Way
41|F775W (HST) AB      | 25.21     |+/-0.06 |mag                 |3.86E+14|  2.99E-07|+/-1.65E-08|Jy|2011ApJ...738...69S|uncertainty|      7764 A         | Broad-band measurement|03 32 29.29 -27 56 19.46 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
42|F775W (HST/ACS) AB  | 25.12     ||mag                 |3.86E+14|  3.24E-07||Jy|2007A&A...461...39F|no uncertainty reported|    7764   A         | Broad-band measurement|03 32 29.29 -27 56 19.4 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data; derived from a fluxin a different band and a color
43|816 nm              | 1.115E-02 |+/-3.128E-03|photons/m^2^/s/nm   |3.67E+14|  6.03E-07|+/-1.69E-07|Jy|2004A&A...421..913W|1 sigma| 816       nm        | Broad-band measurement|033229.289 -275619.36 (J2000)| Flux in fixed aperture|          0          01.5" aperture     |From new raw data
44|857 nm              | 1.773E-02 |+/-6.477E-03|photons/m^2^/s/nm   |3.50E+14|  1.01E-06|+/-3.68E-07|Jy|2004A&A...421..913W|1 sigma| 857       nm        | Broad-band measurement|033229.289 -275619.36 (J2000)| Flux in fixed aperture|          0          01.5" aperture     |From new raw data
45|I                   | 1.524E-02 |+/-4.035E-03|photons/m^2^/s/nm   |3.50E+14|  8.65E-07|+/-2.29E-07|Jy|2004A&A...421..913W|1 sigma| 857       nm        | Broad-band measurement|033229.289 -275619.36 (J2000)| Flux in fixed aperture|          0          01.5" aperture     |From new raw data
46|914 nm              | 1.658E-02 |+/-1.033E-02|photons/m^2^/s/nm   |3.28E+14|  1.00E-06|+/-6.26E-07|Jy|2004A&A...421..913W|1 sigma| 914       nm        | Broad-band measurement|033229.289 -275619.36 (J2000)| Flux in fixed aperture|          0          01.5" aperture     |From new raw data
47|914 nm              | 1.372E-02 |+/-6.452E-03|photons/m^2^/s/nm   |3.28E+14|  8.31E-07|+/-3.91E-07|Jy|2004A&A...421..913W|1 sigma| 914       nm        | Broad-band measurement|033229.289 -275619.36 (J2000)| Flux in fixed aperture|          0          01.5" aperture     |From new raw data
48|F850LP (HST/ACS) AB | 25.05     ||mag                 |3.17E+14|  3.47E-07||Jy|2004ApJ...600L.119C|no uncertainty reported|    9445   A         | Broad-band measurement|03 32 29.29 -27 56 19.3 (J2000)| Total flux|                                        |Averaged from previously published data
49|F850LP (HST) AB     | 24.86     |+/-0.05 |mag                 |3.17E+14|  4.13E-07|+/-1.90E-08|Jy|2010A&A...510A.109R|uncertainty|      9445 A         | Broad-band measurement|03 32 29.29 -27 56 19.5 (J2000)| Flux in fixed aperture|Corrected to 6" circular aperture       |From reprocessed raw data
50|F850LP (HST/ACS) AB | 24.98     ||mag                 |3.17E+14|  3.70E-07||Jy|2006A&A...454..423V|no uncertainty reported|    9445   A         | Broad-band measurement|033229.29 -275619.5 (J2000)| Total flux|                                        |Averaged new and previously published data
51|F850LP (HST/ACS) AB | 24.984    ||mag                 |3.17E+14|  3.68E-07||Jy|2007A&A...461...39F|no uncertainty reported|    9445   A         | Broad-band measurement|03 32 29.29 -27 56 19.4 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
52|F850LP (HST/ACS) AB | 24.88     |+/-0.04 |mag                 |3.17E+14|  4.05E-07|+/-1.49E-08|Jy|2007ApJ...659...84S|uncertainty|    9445   A         | Broad-band measurement|03 32 29.29 -27 56 19.46 (J2000)| Corrected to total flux from single aperture measurement|                                        |From reprocessed raw data; Extinction-corrected for Milky Way
53|F850LP (HST) AB     | 25.0520   || mag                |3.17E+14|  3.46E-07||Jy|2008A&A...478...83V|no uncertainty reported|      9445 A         | Broad-band measurement|033229.29 -275619.5 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data
54|F850LP (HST) AB     | 25.05     |+/-0.06 |mag                 |3.17E+14|  3.47E-07|+/-1.92E-08|Jy|2011ApJ...738...69S|uncertainty|      9445 A         | Broad-band measurement|03 32 29.29 -27 56 19.46 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
55|J (MUSYC)           ||<1.65      | microJy            |2.42E+14||1.65E-06|Jy|2009MNRAS.395.1905C|3 sigma|      1.24 microns   | Broad-band measurement|03 32 29.30 -27 56 19.40 (J2000)| Not reported in paper|Deboosted flux                          |Averaged from previously published data
56|K (MUSYC)           ||<3.20      | microJy            |1.41E+14||3.20E-06|Jy|2009MNRAS.395.1905C|3 sigma|      2.13 microns   | Broad-band measurement|03 32 29.30 -27 56 19.40 (J2000)| Not reported in paper|Deboosted flux                          |Averaged from previously published data
57|3.6 microns IRAC AB | 23.00     |+/-0.08 |mag                 |8.44E+13|  2.29E-06|+/-1.69E-07|Jy|2010A&A...510A.109R|uncertainty|     3.550 microns   | Broad-band measurement|03 32 29.29 -27 56 19.5 (J2000)| Flux in fixed aperture|Corrected to 6" circular aperture       |From reprocessed raw data
59|3.6 microns IRAC AB | 22.64     |+/-0.02 |mag                 |8.44E+13|  3.19E-06|+/-5.88E-08|Jy|2007ApJ...659...84S|uncertainty|   3.550   microns   | Broad-band measurement|03 32 29.29 -27 56 19.46 (J2000)| Corrected to total flux from single aperture measurement|                                        |From reprocessed raw data
60|3.6 microns IRAC AB | 22.56     |+/-0.06 |mag                 |8.44E+13|  3.44E-06|+/-1.90E-07|Jy|2011ApJ...738...69S|uncertainty|     3.550 microns   | Broad-band measurement|03 32 29.29 -27 56 19.46 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
61|3.6 microns (IRAC)  | 2.48      |+/-0.15 | microJy            |8.44E+13|  2.48E-06|+/-1.50E-07|Jy|2008ApJ...680..130C|1 sigma|     3.550 microns   | Broad-band measurement|53.122323 -27.938676 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
62|4.5 microns IRAC AB | 22.55     |+/-0.02 |mag                 |6.67E+13|  3.47E-06|+/-6.39E-08|Jy|2007ApJ...659...84S|uncertainty|   4.493   microns   | Broad-band measurement|03 32 29.29 -27 56 19.46 (J2000)| Corrected to total flux from single aperture measurement|                                        |From reprocessed raw data
64|4.5 microns (IRAC)  | 2.64      |+/-0.14 | microJy            |6.67E+13|  2.64E-06|+/-1.40E-07|Jy|2008ApJ...680..130C|1 sigma|     4.493 microns   | Broad-band measurement|53.122323 -27.938676 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
65|4.5 microns IRAC AB | 23.05     |+/-0.12 |mag                 |6.67E+13|  2.19E-06|+/-2.42E-07|Jy|2010A&A...510A.109R|uncertainty|     4.493 microns   | Broad-band measurement|03 32 29.29 -27 56 19.5 (J2000)| Flux in fixed aperture|Corrected to 6" circular aperture       |From reprocessed raw data
66|4.5 microns IRAC AB | 22.47     |+/-0.06 |mag                 |6.67E+13|  3.73E-06|+/-2.06E-07|Jy|2011ApJ...738...69S|uncertainty|     4.493 microns   | Broad-band measurement|03 32 29.29 -27 56 19.46 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
67|5.8 microns (IRAC)  | 4.13      |+/-0.46 | microJy            |5.23E+13|  4.13E-06|+/-4.60E-07|Jy|2008ApJ...680..130C|1 sigma|     5.731 microns   | Broad-band measurement|53.122323 -27.938676 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
69|5.8 microns IRAC AB | 21.81     |+/-0.09 |mag                 |5.23E+13|  6.86E-06|+/-5.68E-07|Jy|2011ApJ...738...69S|uncertainty|     5.731 microns   | Broad-band measurement|03 32 29.29 -27 56 19.46 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
70|5.8 microns IRAC AB | 22.52     |+/-0.25 |mag                 |5.23E+13|  3.57E-06|+/-8.21E-07|Jy|2010A&A...510A.109R|uncertainty|     5.731 microns   | Broad-band measurement|03 32 29.29 -27 56 19.5 (J2000)| Flux in fixed aperture|Corrected to 6" circular aperture       |From reprocessed raw data
71|8.0 microns (IRAC)  | 6.44      |+/-0.29 | microJy            |3.81E+13|  6.44E-06|+/-2.90E-07|Jy|2008ApJ...680..130C|1 sigma|     7.872 microns   | Broad-band measurement|53.122323 -27.938676 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
72|8.0 microns IRAC AB | 21.31     |+/-0.24 |mag                 |3.81E+13|  1.09E-05|+/-2.40E-06|Jy|2010A&A...510A.109R|uncertainty|     7.872 microns   | Broad-band measurement|03 32 29.29 -27 56 19.5 (J2000)| Flux in fixed aperture|Corrected to 6" circular aperture       |From reprocessed raw data
74|8.0 microns IRAC AB | 21.30     |+/-0.07 |mag                 |3.81E+13|  1.10E-05|+/-7.07E-07|Jy|2011ApJ...738...69S|uncertainty|     7.872 microns   | Broad-band measurement|03 32 29.29 -27 56 19.46 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
75|24 microns (MIPS)   | 31.60     |+/-5.14 | microJy            |1.27E+13|  3.16E-05|+/-5.14E-06|Jy|2008ApJ...680..130C|1 sigma|     23.68 microns   | Broad-band measurement|53.122323 -27.938676 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
76|24 microns (MIPS)   | 35.6      |+/-2.9  |microJy             |1.27E+13|  3.56E-05|+/-2.90E-06|Jy|2011A&A...528A..35M|uncertainty|     23.68 microns   | Broad-band measurement|03 32 29.29 -27 56 19.00 (J2000)| Flux integrated from map|                                        |From new raw data
77|70 microns (MIPS)   ||<2500      | microJy            |4.20E+12||2.50E-03|Jy|2009MNRAS.395.1905C|3 sigma|     71.42 microns   | Broad-band measurement|03 32 29.30 -27 56 19.40 (J2000)| Not reported in paper|Deboosted flux                          |From new raw data
78|70 microns (MIPS)   ||<4.2       |milliJy             |4.20E+12||4.20E-03|Jy|2011A&A...528A..35M|no uncertainty reported|     71.42 microns   | Broad-band measurement|03 32 29.29 -27 56 19.00 (J2000)| Flux integrated from map|                                        |From new raw data
79|160 microns (MIPS)  ||<33000     | microJy            |1.92E+12||3.30E-02|Jy|2009MNRAS.395.1905C|3 sigma|     155.9 microns   | Broad-band measurement|03 32 29.30 -27 56 19.40 (J2000)| Not reported in paper|Deboosted flux                          |From new raw data
80|[C II] 157.74 (APEX)| 14.7      |+/-2.2  |Jy km/s             |1.90E+12|  1.62E+07|+/-2.42E+06|Jy-Hz|2011A&A...530L...8D|uncertainty| 157.74    microns   | Line measurement; flux integrated over line; lines measured in emission|03 32 29.4 -27 56 19 (J2000)| Flux integrated from map|                                        |From new raw data
81|870 microns (LABOCA)| 5.8       |+/-1.3  |milliJy             |3.45E+11|  5.80E-03|+/-1.30E-03|Jy|2009ApJ...707.1201W|uncertainty|       870 microns   | Broad-band measurement|03 32 29.33 -27 56 19.3 (J2000)| Flux integrated from map|S/N = 4.6                               |From new raw data
82|870 microns (APEX)  | 5000      |+/-1400 | microJy            |3.45E+11|  5.00E-03|+/-1.40E-03|Jy|2009MNRAS.395.1905C|uncertainty|       870 microns   | Broad-band measurement|03 32 29.30 -27 56 19.40 (J2000)| Not reported in paper|Deboosted flux                          |From new raw data
83|1.1 mm (ASTE)       | 3.3       |+/-0.5  |milliJy             |2.73E+11|  3.30E-03|+/-5.00E-04|Jy|2011ApJ...730L..28G|uncertainty|     1.1   mm        | Broad-band measurement|03 32 29.29 -27 56 19.5 (J2000)| From fitting to map|                                        |Averaged from previously published data
84|CO(2-1) (ATCA)      | 0.09      |+/-0.02 |Jy km/s             |2.31E+11|  1.20E+04|+/-2.67E+03|Jy-Hz|2010MNRAS.407L.103C|uncertainty|   230.538 GHz       | Line measurement; flux integrated over line; lines measured in emission|03 32 29.30 -27 56 19.40 (J2000)| Flux integrated from map|                                        |From new raw data
85|20 cm (VLA)         | 18.8      |+/-6.3  | microJy            |1.40E+09|  1.88E-05|+/-6.30E-06|Jy|2009MNRAS.395.1905C|uncertainty|        20 cm        | Broad-band measurement|03 32 29.30 -27 56 19.40 (J2000)| Not reported in paper|Deboosted flux                          |From new raw data
