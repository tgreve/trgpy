
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-06-16T05:27:17PDT



Photometric Data for SDSS J141824.67+523255.4

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|u (SDSS PSF) AB     | 24.478    |+/-1.067|asinh mag           |8.36E+14|  1.53E-07|+/-1.05E-06|Jy|2007SDSS6.C...0000:|based on count statistics only|3585       A         | Broad-band measurement|214.6028133943 52.5487352116 (J2000)| Modelled datum|SDSS flags: CANONICAL_CENTER - used canonical, not local, center; CHILD - object is part of a blended parent object; NOPETRO - no Petrosian radius could be determined; MANYR90 - more than one 90% radius; PETROFAINT - Petrosian radius measured at very low surface brightness; ELLIPFAINT - no isophotal fits performed; AMOMENT_FAINT - too faint for adaptive moments;|From new raw data
2|u (SDSS CModel) AB  | 22.450    ||asinh mag           |8.36E+14|  3.87E-06||Jy|2007SDSS6.C...0000:|no uncertainty reported|3585       A         | Broad-band measurement|214.6028133943 52.5487352116 (J2000)| Modelled datum|SDSS flags: CANONICAL_CENTER - used canonical, not local, center; CHILD - object is part of a blended parent object; NOPETRO - no Petrosian radius could be determined; MANYR90 - more than one 90% radius; PETROFAINT - Petrosian radius measured at very low surface brightness; ELLIPFAINT - no isophotal fits performed; AMOMENT_FAINT - too faint for adaptive moments;|From new raw data
3|u (SDSS Model) AB   | 23.939    |+/-1.815|asinh mag           |8.36E+14|  7.23E-07|+/-2.14E-06|Jy|2007SDSS6.C...0000:|based on count statistics only|3585       A         | Broad-band measurement|214.6028133943 52.5487352116 (J2000)| Modelled datum|SDSS flags: CANONICAL_CENTER - used canonical, not local, center; CHILD - object is part of a blended parent object; NOPETRO - no Petrosian radius could be determined; MANYR90 - more than one 90% radius; PETROFAINT - Petrosian radius measured at very low surface brightness; ELLIPFAINT - no isophotal fits performed; AMOMENT_FAINT - too faint for adaptive moments;|From new raw data
4|g (SDSS PSF) AB     | 24.389    |+/-0.580|asinh mag           |6.17E+14|  4.70E-07|+/-4.30E-07|Jy|2007SDSS6.C...0000:|based on count statistics only|4858       A         | Broad-band measurement|214.6028133943 52.5487352116 (J2000)| Modelled datum|SDSS flags: CANONICAL_CENTER - used canonical, not local, center; CHILD - object is part of a blended parent object; NOPETRO - no Petrosian radius could be determined; NOPETRO_BIG - Petrosian radius is larger than extracted radial profile; MANYR50 - more than one 50% radius; ELLIPFAINT - no isophotal fits performed; AMOMENT_FAINT - too faint for adaptive moments;|From new raw data
5|g (SDSS CModel) AB  | 23.994    ||asinh mag           |6.17E+14|  8.01E-07||Jy|2007SDSS6.C...0000:|no uncertainty reported|4858       A         | Broad-band measurement|214.6028133943 52.5487352116 (J2000)| Modelled datum|SDSS flags: CANONICAL_CENTER - used canonical, not local, center; CHILD - object is part of a blended parent object; NOPETRO - no Petrosian radius could be determined; NOPETRO_BIG - Petrosian radius is larger than extracted radial profile; MANYR50 - more than one 50% radius; ELLIPFAINT - no isophotal fits performed; AMOMENT_FAINT - too faint for adaptive moments;|From new raw data
6|g (SDSS Model) AB   | 23.703    |+/-0.806|asinh mag           |6.17E+14|  1.11E-06|+/-9.56E-07|Jy|2007SDSS6.C...0000:|based on count statistics only|4858       A         | Broad-band measurement|214.6028133943 52.5487352116 (J2000)| Modelled datum|SDSS flags: CANONICAL_CENTER - used canonical, not local, center; CHILD - object is part of a blended parent object; NOPETRO - no Petrosian radius could be determined; NOPETRO_BIG - Petrosian radius is larger than extracted radial profile; MANYR50 - more than one 50% radius; ELLIPFAINT - no isophotal fits performed; AMOMENT_FAINT - too faint for adaptive moments;|From new raw data
7|r (SDSS CModel) AB  | 21.936    ||asinh mag           |4.77E+14|  6.07E-06||Jy|2007SDSS6.C...0000:|no uncertainty reported|6290       A         | Broad-band measurement|214.6028133943 52.5487352116 (J2000)| Modelled datum|SDSS flags: CHILD - object is part of a blended parent object; NOPETRO - no Petrosian radius could be determined; PETROFAINT - Petrosian radius measured at very low surface brightness; ELLIPFAINT - no isophotal fits performed; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding; BRIGHTEST_GALAXY_CHILD - brightest child among one parent's children; CANONICAL_BAND - this band was primary (usually r); AMOMENT_FAINT - too faint for adaptive moments;|From new raw data
8|r (SDSS PSF) AB     | 22.910    |+/-0.251|asinh mag           |4.77E+14|  2.41E-06|+/-5.93E-07|Jy|2007SDSS6.C...0000:|based on count statistics only|6290       A         | Broad-band measurement|214.6028133943 52.5487352116 (J2000)| Modelled datum|SDSS flags: CHILD - object is part of a blended parent object; NOPETRO - no Petrosian radius could be determined; PETROFAINT - Petrosian radius measured at very low surface brightness; ELLIPFAINT - no isophotal fits performed; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding; BRIGHTEST_GALAXY_CHILD - brightest child among one parent's children; CANONICAL_BAND - this band was primary (usually r); AMOMENT_FAINT - too faint for adaptive moments;|From new raw data
9|r (SDSS Model) AB   | 21.936    |+/-0.245|asinh mag           |4.77E+14|  6.07E-06|+/-1.38E-06|Jy|2007SDSS6.C...0000:|based on count statistics only|6290       A         | Broad-band measurement|214.6028133943 52.5487352116 (J2000)| Modelled datum|SDSS flags: CHILD - object is part of a blended parent object; NOPETRO - no Petrosian radius could be determined; PETROFAINT - Petrosian radius measured at very low surface brightness; ELLIPFAINT - no isophotal fits performed; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding; BRIGHTEST_GALAXY_CHILD - brightest child among one parent's children; CANONICAL_BAND - this band was primary (usually r); AMOMENT_FAINT - too faint for adaptive moments;|From new raw data
10|i (SDSS PSF) AB     | 24.925    |+/-0.741|asinh mag           |3.89E+14| -7.09E-07|+/-1.01E-06|Jy|2007SDSS6.C...0000:|based on count statistics only|7706       A         | Broad-band measurement|214.6028133943 52.5487352116 (J2000)| Modelled datum|SDSS flags: CANONICAL_CENTER - used canonical, not local, center; CHILD - object is part of a blended parent object; NOPETRO - no Petrosian radius could be determined; INTERP - object contains interpolated-over pixels; PETROFAINT - Petrosian radius measured at very low surface brightness; ELLIPFAINT - no isophotal fits performed; AMOMENT_FAINT - too faint for adaptive moments;|From new raw data
11|i (SDSS CModel) AB  | 24.878    ||asinh mag           |3.89E+14| -6.45E-07||Jy|2007SDSS6.C...0000:|no uncertainty reported|7706       A         | Broad-band measurement|214.6028133943 52.5487352116 (J2000)| Modelled datum|SDSS flags: CANONICAL_CENTER - used canonical, not local, center; CHILD - object is part of a blended parent object; NOPETRO - no Petrosian radius could be determined; INTERP - object contains interpolated-over pixels; PETROFAINT - Petrosian radius measured at very low surface brightness; ELLIPFAINT - no isophotal fits performed; AMOMENT_FAINT - too faint for adaptive moments;|From new raw data
12|i (SDSS Model) AB   | 25.027    |+/-1.512|asinh mag           |3.89E+14| -8.52E-07|+/-2.17E-06|Jy|2007SDSS6.C...0000:|based on count statistics only|7706       A         | Broad-band measurement|214.6028133943 52.5487352116 (J2000)| Modelled datum|SDSS flags: CANONICAL_CENTER - used canonical, not local, center; CHILD - object is part of a blended parent object; NOPETRO - no Petrosian radius could be determined; INTERP - object contains interpolated-over pixels; PETROFAINT - Petrosian radius measured at very low surface brightness; ELLIPFAINT - no isophotal fits performed; AMOMENT_FAINT - too faint for adaptive moments;|From new raw data
13|z (SDSS PSF) AB     | 21.912    |+/-0.493|asinh mag           |3.25E+14|  4.99E-06|+/-3.30E-06|Jy|2007SDSS6.C...0000:|based on count statistics only|9222       A         | Broad-band measurement|214.6028133943 52.5487352116 (J2000)| Modelled datum|SDSS flags: CANONICAL_CENTER - used canonical, not local, center; CHILD - object is part of a blended parent object; ELLIPFAINT - no isophotal fits performed; BINNED1 - detected at >=5 sigma in original imaging frame; DEBLEND_NOPEAK - object has no detected peak;|From new raw data
14|z (SDSS CModel) AB  | 21.999    ||asinh mag           |3.25E+14|  4.42E-06||Jy|2007SDSS6.C...0000:|no uncertainty reported|9222       A         | Broad-band measurement|214.6028133943 52.5487352116 (J2000)| Modelled datum|SDSS flags: CANONICAL_CENTER - used canonical, not local, center; CHILD - object is part of a blended parent object; ELLIPFAINT - no isophotal fits performed; BINNED1 - detected at >=5 sigma in original imaging frame; DEBLEND_NOPEAK - object has no detected peak;|From new raw data
15|z (SDSS Model) AB   | 21.947    |+/-1.240|asinh mag           |3.25E+14|  4.76E-06|+/-8.12E-06|Jy|2007SDSS6.C...0000:|based on count statistics only|9222       A         | Broad-band measurement|214.6028133943 52.5487352116 (J2000)| Modelled datum|SDSS flags: CANONICAL_CENTER - used canonical, not local, center; CHILD - object is part of a blended parent object; ELLIPFAINT - no isophotal fits performed; BINNED1 - detected at >=5 sigma in original imaging frame; DEBLEND_NOPEAK - object has no detected peak;|From new raw data
16|K_s (Keck)          | 18.53     || mag                |1.39E+14|  2.40E-05||Jy|2007MNRAS.382..109T|no uncertainty reported|      2.15 microns   | Broad-band measurement|214.60303 +52.54876 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
17|CO(3-2) (PdBI)      ||<0.06      |Jy km/s             |3.46E+11|  1.52E+05|3.04E+04|Jy-Hz|2010Natur.463..781T|3 sigma|   345.998 GHz       | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|                                        |From new raw data
