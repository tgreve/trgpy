
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-07-10T13:02:05PDT



Photometric Data for LEDA 2831332

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|3.6 microns (IRAC)  | 61.6      |+/-6.4  | microJy            |8.44E+13|  6.16E-05|+/-6.40E-06|Jy|2007ApJS..171..353S|uncertainty|   3.550   microns   | Broad-band measurement|22 27 43.3 -27 05 01.71 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
2|4.5 microns (IRAC)  | 86.1      |+/-8.8  | microJy            |6.67E+13|  8.61E-05|+/-8.80E-06|Jy|2007ApJS..171..353S|uncertainty|   4.493   microns   | Broad-band measurement|22 27 43.3 -27 05 01.71 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
3|5.8 microns (IRAC)  | 98.4      |+/-10.0 | microJy            |5.23E+13|  9.84E-05|+/-1.00E-05|Jy|2007ApJS..171..353S|uncertainty|   5.731   microns   | Broad-band measurement|22 27 43.3 -27 05 01.71 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
4|8.0 microns (IRAC)  | 203.9     |+/-20.5 | microJy            |3.81E+13|  2.04E-04|+/-2.05E-05|Jy|2007ApJS..171..353S|uncertainty|   7.872   microns   | Broad-band measurement|22 27 43.3 -27 05 01.71 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
5|1.4GHz (VLA)        | 269.9     |+/-8.1  |milliJy             |1.40E+09|  2.70E-01|+/-8.10E-03|Jy|1998AJ....115.1693C|uncertainty|    1.40   GHz       | Broad-band measurement|22 27 43.26 -27 05 1.3 (J2000)| Flux integrated from map|                                        |From new raw data
6|408 MHz             | 1.15      |+/-0.07 |Jy                  |4.08E+08|  1.15E+00|+/-7.00E-02|Jy|1981MNRAS.194..693L|rms noise|408        MHz       | Broad-band measurement|222455.9 -272034 (B1950)| Modelled datum|                                        |From new raw data; Corrected for contaminating sources
7|365 MHz (Texas)     | 1.092     |+/-0.032|Jy                  |3.65E+08|  1.09E+00|+/-3.20E-02|Jy|1996AJ....111.1945D|internal error|365        MHz       | Broad-band measurement; obtained by interpolation over frequency|222455.893 -272022.43 (B1950)| Integrated from scans|Model:P;MFlag:+;EFlag:+;LFlag:+.        |From new raw data
8|74 MHz (VLA)        | 0.61      |+/-0.10 | Jy                 |7.38E+07|  6.10E-01|+/-1.00E-01|Jy|2007AJ....134.1245C|rms uncertainty|      73.8 MHz       | Broad-band measurement|22 27 43.18 -27 05 00.8 (J2000)| Flux integrated from map|Corrected for clean bias                |From new raw data
