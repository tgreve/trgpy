
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-07-08T07:37:11PDT



Photometric Data for LBQS 0018-0220

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|Photographic IIIa-J | 17.44     |+/-0.15 |mag                 |6.48E+14|  4.50E-04|+/-6.67E-05|Jy|1995AJ....109.1498H|estimated error|4627       A         | Broad-band measurement; photometric system transformed|001853.83 -022012.1 (B1950)| Integrated from scans|                                        |From new raw data; Uncorrected for known sources in beam
4|350 microns (CSO/SHARC)   | 32        |+/-5    |milliJy             |8.57E+11|  3.20E-02|+/-5.00E-03|Jy|2009ApJ...707..988W|rms noise|       350 microns   | Broad-band measurement|00 21 27.30 -02 03 33.0 (J2000)| Flux integrated from map|S/N=6.4 sigma                           |From new raw data
5|350 GHz 850um (SCUBA)     | 17.2      |+/-2.9  |milliJy             |3.50E+11|  1.72E-02|+/-2.90E-03|Jy|2006AJ....132.1307P|uncertainty|     350   GHz       | Broad-band measurement|00 21 27.37 -02 03 33.8 (J2000)| Flux integrated from map|From 2003MNRAS.339.1183P                |Averaged from previously published data; OBJ_NAME modifiedfrom published value
7|5.0 GHz (VLA)       ||<120E-06   |Jy                  |5.00E+09||1.20E-04|Jy|2006AJ....132.1307P|3 sigma|     5.0   GHz       | Broad-band measurement|00 21 27.37 -02 03 33.8 (J2000)| Flux integrated from map|                                        |From new raw data; OBJ_NAME modified from published value
8|1.4 GHz (VLA)       | 260E-06   |+/-20E-06|Jy                  |1.40E+09|  2.60E-04|+/-2.00E-05|Jy|2006AJ....132.1307P|1 sigma|     1.4   GHz       | Broad-band measurement|00 21 27.37 -02 03 33.8 (J2000)| Flux integrated from map|                                        |From new raw data; OBJ_NAME modified from published value
