
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-07-08T05:16:52PDT



Photometric Data for GOODS J123721.45+621346.5

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|NUV (GALEX) AB      | 24.53     |+/-0.10 |mag                 |1.95E+15|  5.60E-07|+/-5.16E-08|Jy|2011ApJ...734L..12B|uncertainty|      1539 A         | Broad-band measurement|12 37 21.4 +62 13 46.1 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
2|U (KPNO) AB         | 24.41     |+/-0.11 |mag                 |8.44E+14|  6.25E-07|+/-6.33E-08|Jy|2011ApJ...734L..12B|uncertainty|      3552 A         | Broad-band measurement|12 37 21.4 +62 13 46.1 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
3|U (KPNO) AB         | 24.5      || mag                |8.22E+14|  5.76E-07||Jy|2004AJ....127.3137C|no uncertainty reported| 3647.65   A         | Broad-band measurement|189.339386 +62.22958 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
4|B (HST/ACS) AB      | 24.336    ||mag                 |6.98E+14|  6.69E-07||Jy|2007ApJ...660...81M|no uncertainty reported|    4297   A         | Broad-band measurement|12 37 21.474 +62 13 46.03 (J2000)| Flux integrated from map|                                        |From reprocessed raw data; Corrected for contaminatingsources
5|B (Subaru) AB       | 24.5      || mag                |6.77E+14|  5.76E-07||Jy|2004AJ....127.3137C|no uncertainty reported| 4427.60   A         | Broad-band measurement|189.339386 +62.22958 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
6|B (Subaru) AB       | 24.47     ||mag                 |6.77E+14|  5.92E-07||Jy|2006ApJ...653.1027W|no uncertainty reported| 4427.60   A         | Broad-band measurement|189.339475 62.229453 (J2000)| Flux in fixed aperture|3" diameter aperture                    |Averaged from previously published data
7|V (Subaru) AB       | 24.1      || mag                |5.48E+14|  8.32E-07||Jy|2004AJ....127.3137C|no uncertainty reported| 5471.22   A         | Broad-band measurement|189.339386 +62.22958 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
8|V (HST/ACS) AB      | 23.642    ||mag                 |5.08E+14|  1.27E-06||Jy|2007ApJ...660...81M|no uncertainty reported|    5907   A         | Broad-band measurement|12 37 21.474 +62 13 46.03 (J2000)| Flux integrated from map|                                        |From reprocessed raw data; Corrected for contaminatingsources
9|R (Keck II) AB      | 23.72     || mag                |4.62E+14|  1.18E-06||Jy|2004AJ....127.3121W|no uncertainty reported|   648.7   A         | Broad-band measurement|12 37 21.474 +62 13 46.03 (J2000)| Total flux|                                        |From new raw data
10|R (Subaru) AB       | 23.6      || mag                |4.59E+14|  1.32E-06||Jy|2004AJ....127.3137C|no uncertainty reported| 6534.16   A         | Broad-band measurement|189.339386 +62.22958 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
11|R (Subaru) AB       | 23.58     ||mag                 |4.59E+14|  1.34E-06||Jy|2006ApJ...653.1027W|no uncertainty reported| 6534.16   A         | Broad-band measurement|189.339475 62.229453 (J2000)| Flux in fixed aperture|3" diameter aperture                    |Averaged from previously published data
12|i (HST/ACS) AB      | 22.702    ||mag                 |3.86E+14|  3.01E-06||Jy|2007ApJ...660...81M|no uncertainty reported|    7764   A         | Broad-band measurement|12 37 21.474 +62 13 46.03 (J2000)| Flux integrated from map|                                        |From reprocessed raw data; Corrected for contaminatingsources
13|I (Subaru) AB       | 22.7      || mag                |3.76E+14|  3.02E-06||Jy|2004AJ....127.3137C|no uncertainty reported| 7975.89   A         | Broad-band measurement|189.339386 +62.22958 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
14|I (Subaru) AB       | 22.72     ||mag                 |3.76E+14|  2.96E-06||Jy|2006ApJ...653.1027W|no uncertainty reported| 7975.89   A         | Broad-band measurement|189.339475 62.229453 (J2000)| Flux in fixed aperture|3" diameter aperture                    |Averaged from previously published data
15|z' (Subaru) AB      | 22.3      || mag                |3.31E+14|  4.37E-06||Jy|2004AJ....127.3137C|no uncertainty reported| 9069.21   A         | Broad-band measurement|189.339386 +62.22958 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
16|z (HST/ACS) AB      | 22.061    ||mag                 |3.17E+14|  5.44E-06||Jy|2007ApJ...660...81M|no uncertainty reported|    9445   A         | Broad-band measurement|12 37 21.474 +62 13 46.03 (J2000)| Flux integrated from map|                                        |From reprocessed raw data; Corrected for contaminatingsources
17|HK' (UH) AB         | 20.9      || mag                |1.58E+14|  1.59E-05||Jy|2004AJ....127.3137C|no uncertainty reported|18947.38   A         | Broad-band measurement|189.339386 +62.22958 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
18|HK' (QUIRC) AB      | 20.93     |+/-0.12 |mag                 |1.58E+14|  1.54E-05|+/-1.70E-06|Jy|2006ApJ...653.1027W|uncertainty|18947.38   A         | Broad-band measurement|189.339475 62.229453 (J2000)| Flux in fixed aperture|3" diameter aperture                    |Averaged from previously published data
19|3.6 microns (IRAC)  | 45.60     |+/-2.28 |microJy             |8.44E+13|  4.56E-05|+/-2.28E-06|Jy|2011AJ....141....1T|rms uncertainty|     3.550 microns   | Broad-band measurement|189.339371 62.229511 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
20|4.5 microns (IRAC)  | 36.20     |+/-1.81 |microJy             |6.67E+13|  3.62E-05|+/-1.81E-06|Jy|2011AJ....141....1T|rms uncertainty|     4.493 microns   | Broad-band measurement|189.339371 62.229511 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
21|5.8 microns (IRAC)  | 27.10     |+/-1.40 |microJy             |5.23E+13|  2.71E-05|+/-1.40E-06|Jy|2011AJ....141....1T|rms uncertainty|     5.731 microns   | Broad-band measurement|189.339371 62.229511 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
22|8.0 microns (IRAC)  | 27.00     |+/-1.42 |microJy             |3.81E+13|  2.70E-05|+/-1.42E-06|Jy|2011AJ....141....1T|rms uncertainty|     7.872 microns   | Broad-band measurement|189.339371 62.229511 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
23|16 microns (IRS)    | 212.1     |+/-9.1  |microJy             |1.90E+13|  2.12E-04|+/-9.10E-06|Jy|2011AJ....141....1T|rms uncertainty|      15.8 microns   | Broad-band measurement|189.339371 62.229511 (J2000)| From fitting to map|                                        |From new raw data
24|24 microns (MIPS)   | 235.0     |+/-7.5  |microJy             |1.27E+13|  2.35E-04|+/-7.50E-06|Jy|2011AJ....141....1T|rms uncertainty|     23.68 microns   | Broad-band measurement|189.339371 62.229511 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
25|24 microns (MIPS)   | 217       |+/-6    |microJy             |1.27E+13|  2.17E-04|+/-6.00E-06|Jy|2011ApJ...726...93R|uncertainty|     23.68 microns   | Broad-band measurement|12 37 21.45 +62 13 46.1 (J2000)| Not reported in paper|                                        |Averaged from previously published data
26|24 microns (MIPS)   | 235.0     |+/-7.5  |microJy             |1.27E+13|  2.35E-04|+/-7.50E-06|Jy|2011ApJ...734L..12B|uncertainty|     23.68 microns   | Broad-band measurement|12 37 21.4 +62 13 46.1 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
27|24 microns (MIPS)   | 239.5     |+/-4.2  |microJy             |1.27E+13|  2.40E-04|+/-4.20E-06|Jy|2011A&A...528A..35M|uncertainty|     23.68 microns   | Broad-band measurement|12 37 21.45 +62 13 46.17 (J2000)| Flux integrated from map|                                        |From new raw data
1|MIPS 24 microns      | 238.    |+/-8.0 |microJy         |1.25E+13 |  238.E-06|+/-8.0E-06 |Jy|1990IRASF.C...0000M|3sigma uncertainty| 25        microns   | Broad-band measurement|115813.1 +302058 (B1950)| Flux in fixed aperture|                                        |From new raw data
28|70 microns (MIPS)   ||<5.8       |milliJy             |4.20E+12||5.80E-03|Jy|2011A&A...528A..35M|no uncertainty reported|     71.42 microns   | Broad-band measurement|12 37 21.45 +62 13 46.17 (J2000)| Flux integrated from map|                                        |From new raw data
2|70 microns (PACS)    | 1.8     |+/-0.6 |mJy             |4.283e+12|  1.8E-03 |+/-0.6E-03 |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
3|100 microns (PACS)   | 3.1     |+/-0.3 |mJy             |2.998e+12|  3.1E-03 |+/-0.3E-03 |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
4|160 microns (PACS)   | 8.5     |+/-0.8 |mJy             |1.874e+12|  8.5E-03 |+/-0.8E-03 |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
29|250 microns (SPIRE) | 15.4      |+/-2.6  |milliJy             |1.20E+12|  1.54E-02|+/-2.60E-03|Jy|2011ApJ...734L..12B|uncertainty|       250 microns   | Broad-band measurement|12 37 21.4 +62 13 46.1 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
5|250 microns (SPIRE)  | 14.5    |+/-2.5 |mJy             |1.199e+12|  14.5E-03|+/-2.5e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
6|350 microns (SPIRE)  | 10.8    |+/-3.0 |mJy             |8.565e+11|  10.8E-03|+/-3.0e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
7|500 microns (SPIRE)  | 8.0     |+/-5.0 |mJy             |5.996e+11|  8.0E-03 |5.0e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
8|1160 microns (Penner)|         |<1.6   |mJy             |2.58442e+08|        |1.6E-03|Jy |2.40e+01 |3sigma |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
8|1160 microns (Penner)|         |<1.6   |mJy             |2.58442E+11|       |1.6E-03|Jy|2004MNRAS.354..779G|3sigma uncertainty|      1200 microns   | Broad-band measurement|16 36 55.9 +40 59 12 (J2000)| Flux integrated from map|S/N = 3.66                              |From new raw data
30|1.4 GHz (VLA)       | 41.6      |+/-8.7  |microJy             |1.40E+09|  4.16E-05|+/-8.70E-06|Jy|2010ApJS..188..178M|uncertainty|       1.4 GHz       | Broad-band measurement|12 37 21.45 +62 13 46.1 (J2000)| Total flux; Beam filling or dilution corrected|Major=1.0"; Minor=0.1"; PA=27 deg       |From new raw data
31|1.4 GHz (VLA)       | 50        ||microJy             |1.40E+09|  5.00E-05||Jy|2005MNRAS.358.1159M|no uncertainty reported|     1.4   GHz       | Broad-band measurement|12 37 21.4669 +62 13 46.675 (J2000)| Flux integrated from map|                                        |From new raw data
32|1.4 GHz (VLA)       | 47        |+/-12   | microJy            |1.40E+09|  4.70E-05|+/-1.20E-05|Jy|2006MNRAS.371..963B|1 sigma|       1.4 GHz       | Broad-band measurement|12 37 21.454 +62 13 46.59 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
33|1.4 GHz (VLA)       | 50.5      |+/-8.2  |microJy             |1.40E+09|  5.05E-05|+/-8.20E-06|Jy|2000ApJ...533..611R|1 sigma|1.4        GHz       | Broad-band measurement; broad-band flux derived by integration over spectrum; synthetic band|123721.452 +621346.51 (J2000)| Flux integrated from map; Pointing and beam filling|                                        |From new raw data; Corrected for contaminating sources
