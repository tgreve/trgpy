
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-07-10T13:05:38PDT



Photometric Data for 4C +72.26

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|F702W (HST)         | 8.18      |+/-0.16 |microJy             |4.33E+14|  8.18E-06|+/-1.60E-07|Jy|2010MNRAS.404.1089S|1 sigma|      6919 A         | Broad-band measurement|| Flux in fixed aperture|                                        |From reprocessed raw data
2|K' (Subaru)         | 134       |+/-7    |microJy             |1.41E+14|  1.34E-04|+/-7.00E-06|Jy|2010MNRAS.404.1089S|1 sigma|      2.13 microns   | Broad-band measurement|| Flux in fixed aperture|                                        |From new raw data
3|3.6 microns (IRAC)  | 200.0     |+/-20.0 | microJy            |8.44E+13|  2.00E-04|+/-2.00E-05|Jy|2007ApJS..171..353S|uncertainty|   3.550   microns   | Broad-band measurement|19 08 23.7 +72 20 11.82 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
4|4.5 microns (IRAC)  | 229.0     |+/-23.0 | microJy            |6.67E+13|  2.29E-04|+/-2.30E-05|Jy|2007ApJS..171..353S|uncertainty|   4.493   microns   | Broad-band measurement|19 08 23.7 +72 20 11.82 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
5|5.8 microns (IRAC)  | 241.0     |+/-25.0 | microJy            |5.23E+13|  2.41E-04|+/-2.50E-05|Jy|2007ApJS..171..353S|uncertainty|   5.731   microns   | Broad-band measurement|19 08 23.7 +72 20 11.82 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
6|8.0 microns (IRAC)  | 480.0     |+/-48.0 | microJy            |3.81E+13|  4.80E-04|+/-4.80E-05|Jy|2007ApJS..171..353S|uncertainty|   7.872   microns   | Broad-band measurement|19 08 23.7 +72 20 11.82 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
7|12 microns (ISOCAM) | 0.7       |+/-0.08 |milliJy             |2.50E+13|  7.00E-04|+/-8.00E-05|Jy|2004A&A...421..129S|1 sigma|    12.0   microns   | Broad-band measurement|| From multi-aperture data|                                        |From reprocessed raw data
8|16 microns (IRS)    | 841.0     |+/-70.6 | microJy            |1.87E+13|  8.41E-04|+/-7.06E-05|Jy|2007ApJS..171..353S|uncertainty|      16   microns   | Broad-band measurement|19 08 23.7 +72 20 11.82 (J2000)| Flux in fixed aperture|6" diameter aperture                    |From reprocessed raw data
9|16 microns (IRS)    | 1320      |+/-70   |microJy             |1.87E+13|  1.32E-03|+/-7.00E-05|Jy|2008ApJ...681L...1S|uncertainty|      16   microns   | Broad-band measurement|| Not reported in paper|                                        |From new raw data
10|24 microns (MIPS)   | 1910.0    |+/-98.9 | microJy            |1.27E+13|  1.91E-03|+/-9.89E-05|Jy|2007ApJS..171..353S|uncertainty|   23.68   microns   | Broad-band measurement|19 08 23.7 +72 20 11.82 (J2000)| Flux in fixed aperture|13" diameter aperture                   |From reprocessed raw data
11|70 microns (MIPS)   | 16200     |+/-1905 | microJy            |4.20E+12|  1.62E-02|+/-1.91E-03|Jy|2007ApJS..171..353S|uncertainty|   71.42   microns   | Broad-band measurement|19 08 23.7 +72 20 11.82 (J2000)| Flux in fixed aperture|35" diameter aperture                   |From reprocessed raw data
12|160 microns (MIPS)  ||<63300     | microJy            |1.92E+12||6.33E-02|Jy|2007ApJS..171..353S|3 sigma|   155.9   microns   | Broad-band measurement|19 08 23.7 +72 20 11.82 (J2000)| Flux in fixed aperture|50" diameter aperture                   |From reprocessed raw data
5|250 microns (SPIRE)| 57.2      |+/-2.7 |mJy             |1.199e+12| 57.2E-03|+/-2.7e-03 |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
6|350 microns (SPIRE)| 69.6     |+/-2.8  |mJy             |8.565e+11|69.6E-03 |+/-2.8e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
13|450 microns (SCUBA) | 33        |+/-17   | milliJy            |6.66E+11|  3.30E-02|+/-1.70E-02|Jy|2004MNRAS.353..377R|uncertainty|       450 microns   | Broad-band measurement|19 08 23.70 +72 20 11.8 (J2000)| Not reported in paper|Good quality data                       |From new raw data
8|500 microns (SPIRE) | 63.4     |+/-3.3 |mJy             |5.996e+11|63.4E-03 |+/-3.3e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
14|850 microns (SCUBA) | 10.8      |+/-1.2  | milliJy            |3.53E+11|  1.08E-02|+/-1.20E-03|Jy|2004MNRAS.353..377R|uncertainty|       850 microns   | Broad-band measurement|19 08 23.70 +72 20 11.8 (J2000)| Not reported in paper|Good quality data                       |From new raw data
14|850 microns (SCUBA) | 34.9      |+/-3.0  | milliJy            |3.53E+11|  34.9E-03|+/-3.0E-03|Jy|2004MNRAS.353..377R|uncertainty|       850 microns   | Broad-band measurement|19 08 23.70 +72 20 11.8 (J2000)| Not reported in paper|Good quality data                       |From new raw data
15|4.85 GHz            | 53        |+/-6    |milliJy             |4.85E+09|  5.30E-02|+/-6.00E-03|Jy|1991ApJS...75.1011G|rms noise|4.85       GHz       | Broad-band measurement|190907.0 +721515 (B1950)| Modelled datum|                                        |From new raw data; Corrected for contaminating sources
16|4.85 GHz            | 50        |+/-15  %|milliJy             |4.85E+09|  5.00E-02|+/-7.50E-03|Jy|1991ApJS...75....1B|uncertainty|4.85       GHz       | Broad-band measurement|190907.8 +721519 (B1950)| Peak flux|                                        |From new raw data; Corrected for contaminating sources
17|1.40 GHz            | 259       ||milliJy             |1.40E+09|  2.59E-01||Jy|1992ApJS...79..331W|no uncertainty reported|1.4        GHz       | Broad-band measurement|190907.8 +721519 (B1950)| Peak flux|                                        |From new raw data
18|1.4GHz (VLA)        | 296.7     |+/-10.5 |milliJy             |1.40E+09|  2.97E-01|+/-1.05E-02|Jy|1998AJ....115.1693C|uncertainty|    1.40   GHz       | Broad-band measurement|19 08 23.51 +72 20 9.8 (J2000)| Flux integrated from map|                                        |From new raw data
19|92 cm (WENSS)       | 1882      |+/-75.5 |milliJy             |3.25E+08|  1.88E+00|+/-7.55E-02|Jy|1997A&AS..124..259R|uncertainty|92         cm        | Broad-band measurement|190909.42 +721514.2 (B1950)| Flux integrated from map|Single component source                 |From new raw data
20|92 cm (WENSS)       | 1871      |+/-75.1 |milliJy             |3.25E+08|  1.87E+00|+/-7.51E-02|Jy|1997A&AS..124..259R|uncertainty|92         cm        | Broad-band measurement|190909.42 +721514.2 (B1950)| Peak flux|Single component source                 |From new raw data
21|325 MHz (WSRT)      | 1882      || milliJy            |3.25E+08|  1.88E+00||Jy|1997A&AS..124..259R|no uncertainty reported|   325.125 MHz       | Broad-band measurement|19 09 09.42 +72 15 14.2 (B1950)| Flux integrated from map|a=0"; b=0"; PA=0 deg                    |From new raw data
22|178 MHz             | 3.2       |+/-15.0%|Jy                  |1.78E+08|  3.20E+00|+/-4.80E-01|Jy|1967MmRAS..71...49G|uncertainty|178        MHz       | Broad-band measurement|190911.3 +721418 (B1950)| Integrated from scans|                                        |From new raw data; Uncorrected for known sources in beam
23|151 MHz (6C)        | 4.19      |+/-0.040|Jy                  |1.52E+08|  4.19E+00|+/-4.00E-02|Jy|1991MNRAS.251...46H|typical accuracy|151.5      MHz       | Broad-band measurement|190910.1 721514. (B1950)| Peak flux|                                        |From new raw data
24|151 MHz (6C)        | 4.07      |+/-0.090|Jy                  |1.52E+08|  4.07E+00|+/-9.00E-02|Jy|1991MNRAS.251...46H|typical accuracy|151.5      MHz       | Broad-band measurement|190910.1 721514. (B1950)| Flux integrated from map|                                        |From new raw data
25|74 MHz (VLA)        | 8.15      |+/-0.82 | Jy                 |7.38E+07|  8.15E+00|+/-8.20E-01|Jy|2007AJ....134.1245C|rms uncertainty|      73.8 MHz       | Broad-band measurement|19 08 24.29 +72 20 08.9 (J2000)| Flux integrated from map|Corrected for clean bias                |From new raw data
26|38 MHz (8C)         | 11.7      |+/-10.0%|Jy                  |3.78E+07|  1.17E+01|+/-1.17E+00|Jy|1995MNRAS.274..447H|no uncertainty reported|38         MHz       | Broad-band measurement|190909. +721518. (B1950)| Peak flux|Part of multiple component source       |From new raw data
27|38 MHz (8C)         | 14.3      |+/-10.0%|Jy                  |3.78E+07|  1.43E+01|+/-1.43E+00|Jy|1995MNRAS.274..447H|no uncertainty reported|38         MHz       | Broad-band measurement|190909. +721518. (B1950)| Flux integrated from map|Part of multiple component source       |From new raw data
