
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-06-17T09:40:16PDT



Photometric Data for SDF J132415.7+273058

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
2|i' (Subaru) AB      | 27.33     ||mag                 |3.89E+14|  4.25E-08||Jy|2005PASJ...57..165T|no uncertainty reported|    7709   A         | Broad-band measurement|132415.7 +273058 (J2000)| Flux in fixed aperture|2.0" diam aperture                      |From new raw data
3|z' (Subaru) AB      | 25.69     ||mag                 |3.31E+14|  1.92E-07||Jy|2005PASJ...57..165T|no uncertainty reported|    9054   A         | Broad-band measurement|132415.7 +273058 (J2000)| Flux in fixed aperture|2.0" diam aperture                      |From new raw data
4|NB921 (Subaru) AB   | 24.13     ||mag                 |3.26E+14|  8.09E-07||Jy|2005PASJ...57..165T|no uncertainty reported|    9196   A         | Broad-band measurement|132415.7 +273058 (J2000)| Flux in fixed aperture|2.0" diam aperture                      |From new raw data
5|9500 A (Subaru) AB  | 24.73     ||mag                 |3.16E+14|  4.66E-07||Jy|2005PASJ...57..165T|no uncertainty reported|    9500   A         | Broad-band measurement|132415.7 +273058 (J2000)| Flux in fixed aperture|2.0" diam aperture                      |From new raw data; Corrected for flux in reference beam
6|450 microns (SCUBA) | 11.9      ||milliJy             |6.66E+11|  1.19E-02||Jy|2007ApJ...659...76W|no uncertainty reported|     450   microns   | Broad-band measurement|13 24 17.80 +27 30 41.5 (J2000)| Flux integrated from map|S/N = 2.8                               |From new raw data
7|450 microns (SCUBA) ||<9.0       |milliJy             |6.66E+11||9.00E-03|Jy|2007ApJ...659...76W|3 sigma|     450   microns   | Broad-band measurement|13 24 15.7 +27 30 58 (J2000)| Flux integrated from map|                                        |From new raw data
8|850 microns (SCUBA) ||<1.5       |milliJy             |3.53E+11||1.50E-03|Jy|2007ApJ...659...76W|3 sigma|     850   microns   | Broad-band measurement|13 24 15.7 +27 30 58 (J2000)| Flux integrated from map|                                        |From new raw data
9|850 microns (SCUBA) | 5.1       ||milliJy             |3.53E+11|  5.10E-03||Jy|2007ApJ...659...76W|no uncertainty reported|     850   microns   | Broad-band measurement|13 24 17.80 +27 30 41.5 (J2000)| Flux integrated from map|S/N = 7.4                               |From new raw data
11|CARMA 252GHz      |      |<0.37 |mJy                 |2.52E+11|  |0.37E-03|Jy|2011ApJ...736L..28C|1sigma uncertainty|     13006 A         | Broad-band measurement|| Flux in fixed aperture|                                        |From new raw data
