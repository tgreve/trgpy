
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-06-16T16:25:00PDT



Photometric Data for SDSS J142012.98+525613.4

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|u (SDSS PSF) AB     | 22.370    |+/-0.334|asinh mag           |8.36E+14|  4.18E-06|+/-1.33E-06|Jy|2007SDSS6.C...0000:|based on count statistics only|3585       A         | Broad-band measurement|215.0540837723 52.9370608868 (J2000)| Modelled datum|SDSS flags: CANONICAL_CENTER - used canonical, not local, center; NOPETRO - no Petrosian radius could be determined; PETROFAINT - Petrosian radius measured at very low surface brightness; ELLIPFAINT - no isophotal fits performed;|From new raw data
2|u (SDSS CModel) AB  | 22.451    ||asinh mag           |8.36E+14|  3.87E-06||Jy|2007SDSS6.C...0000:|no uncertainty reported|3585       A         | Broad-band measurement|215.0540837723 52.9370608868 (J2000)| Modelled datum|SDSS flags: CANONICAL_CENTER - used canonical, not local, center; NOPETRO - no Petrosian radius could be determined; PETROFAINT - Petrosian radius measured at very low surface brightness; ELLIPFAINT - no isophotal fits performed;|From new raw data
3|u (SDSS Model) AB   | 22.401    |+/-0.415|asinh mag           |8.36E+14|  4.06E-06|+/-1.60E-06|Jy|2007SDSS6.C...0000:|based on count statistics only|3585       A         | Broad-band measurement|215.0540837723 52.9370608868 (J2000)| Modelled datum|SDSS flags: CANONICAL_CENTER - used canonical, not local, center; NOPETRO - no Petrosian radius could be determined; PETROFAINT - Petrosian radius measured at very low surface brightness; ELLIPFAINT - no isophotal fits performed;|From new raw data
4|g (SDSS PSF) AB     | 22.868    |+/-0.128|asinh mag           |6.17E+14|  2.55E-06|+/-3.10E-07|Jy|2007SDSS6.C...0000:|based on count statistics only|4858       A         | Broad-band measurement|215.0540837723 52.9370608868 (J2000)| Modelled datum|SDSS flags: NOPETRO - no Petrosian radius could be determined; PETROFAINT - Petrosian radius measured at very low surface brightness; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
5|g (SDSS CModel) AB  | 21.583    ||asinh mag           |6.17E+14|  8.44E-06||Jy|2007SDSS6.C...0000:|no uncertainty reported|4858       A         | Broad-band measurement|215.0540837723 52.9370608868 (J2000)| Modelled datum|SDSS flags: NOPETRO - no Petrosian radius could be determined; PETROFAINT - Petrosian radius measured at very low surface brightness; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
6|g (SDSS Model) AB   | 22.536    |+/-0.125|asinh mag           |6.17E+14|  3.48E-06|+/-4.08E-07|Jy|2007SDSS6.C...0000:|based on count statistics only|4858       A         | Broad-band measurement|215.0540837723 52.9370608868 (J2000)| Modelled datum|SDSS flags: NOPETRO - no Petrosian radius could be determined; PETROFAINT - Petrosian radius measured at very low surface brightness; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
7|r (SDSS CModel) AB  | 22.119    ||asinh mag           |4.77E+14|  5.12E-06||Jy|2007SDSS6.C...0000:|no uncertainty reported|6290       A         | Broad-band measurement|215.0540837723 52.9370608868 (J2000)| Modelled datum|SDSS flags: BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding; CANONICAL_BAND - this band was primary (usually r);|From new raw data
8|r (SDSS PSF) AB     | 22.390    |+/-0.144|asinh mag           |4.77E+14|  3.97E-06|+/-5.39E-07|Jy|2007SDSS6.C...0000:|based on count statistics only|6290       A         | Broad-band measurement|215.0540837723 52.9370608868 (J2000)| Modelled datum|SDSS flags: BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding; CANONICAL_BAND - this band was primary (usually r);|From new raw data
9|r (SDSS Model) AB   | 22.119    |+/-0.146|asinh mag           |4.77E+14|  5.12E-06|+/-6.98E-07|Jy|2007SDSS6.C...0000:|based on count statistics only|6290       A         | Broad-band measurement|215.0540837723 52.9370608868 (J2000)| Modelled datum|SDSS flags: BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding; CANONICAL_BAND - this band was primary (usually r);|From new raw data
10|i (SDSS PSF) AB     | 22.095    |+/-0.169|asinh mag           |3.89E+14|  5.19E-06|+/-8.33E-07|Jy|2007SDSS6.C...0000:|based on count statistics only|7706       A         | Broad-band measurement|215.0540837723 52.9370608868 (J2000)| Modelled datum|SDSS flags: ELLIPFAINT - no isophotal fits performed; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
11|i (SDSS CModel) AB  | 21.739    ||asinh mag           |3.89E+14|  7.26E-06||Jy|2007SDSS6.C...0000:|no uncertainty reported|7706       A         | Broad-band measurement|215.0540837723 52.9370608868 (J2000)| Modelled datum|SDSS flags: ELLIPFAINT - no isophotal fits performed; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
12|i (SDSS Model) AB   | 21.839    |+/-0.175|asinh mag           |3.89E+14|  6.61E-06|+/-1.09E-06|Jy|2007SDSS6.C...0000:|based on count statistics only|7706       A         | Broad-band measurement|215.0540837723 52.9370608868 (J2000)| Modelled datum|SDSS flags: ELLIPFAINT - no isophotal fits performed; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
13|z (SDSS PSF) AB     | 21.630    |+/-0.408|asinh mag           |3.25E+14|  7.07E-06|+/-3.31E-06|Jy|2007SDSS6.C...0000:|based on count statistics only|9222       A         | Broad-band measurement|215.0540837723 52.9370608868 (J2000)| Modelled datum|SDSS flags: CANONICAL_CENTER - used canonical, not local, center; ELLIPFAINT - no isophotal fits performed; AMOMENT_SHIFT - center moved too far while determining adaptive moments;|From new raw data
14|z (SDSS CModel) AB  | 19.204    ||asinh mag           |3.25E+14|  7.41E-05||Jy|2007SDSS6.C...0000:|no uncertainty reported|9222       A         | Broad-band measurement|215.0540837723 52.9370608868 (J2000)| Modelled datum|SDSS flags: CANONICAL_CENTER - used canonical, not local, center; ELLIPFAINT - no isophotal fits performed; AMOMENT_SHIFT - center moved too far while determining adaptive moments;|From new raw data
15|z (SDSS Model) AB   | 21.071    |+/-0.343|asinh mag           |3.25E+14|  1.28E-05|+/-4.37E-06|Jy|2007SDSS6.C...0000:|based on count statistics only|9222       A         | Broad-band measurement|215.0540837723 52.9370608868 (J2000)| Modelled datum|SDSS flags: CANONICAL_CENTER - used canonical, not local, center; ELLIPFAINT - no isophotal fits performed; AMOMENT_SHIFT - center moved too far while determining adaptive moments;|From new raw data
