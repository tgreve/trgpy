
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-06-11T20:42:09PDT



Photometric Data for BzK25536 (z=1.459)

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|R (Keck II) AB      | 25.29     | | mag                |4.62E+14|  2.78E-07| |Jy|2004AJ....127.3121W|no uncertainty reported|   648.7   A         | Broad-band measurement|12 37 28.313 +62 18 54.58 (J2000)| Total flux|                                        |From new raw data
2|3.6 microns (IRAC)  | 22.20     |+/-1.11 |microJy             |8.44E+13|  2.22E-05|+/-1.11E-06|Jy|2011AJ....141....1T|rms uncertainty|     3.550 microns   | Broad-band measurement|189.367981 62.315258 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
3|4.5 microns (IRAC)  | 23.70     |+/-1.19 |microJy             |6.67E+13|  2.37E-05|+/-1.19E-06|Jy|2011AJ....141....1T|rms uncertainty|     4.493 microns   | Broad-band measurement|189.367981 62.315258 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
4|5.8 microns (IRAC)  | 18.00     |+/-1.00 |microJy             |5.23E+13|  1.80E-05|+/-1.00E-06|Jy|2011AJ....141....1T|rms uncertainty|     5.731 microns   | Broad-band measurement|189.367981 62.315258 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
5|8.0 microns (IRAC)  | 14.60     |+/-0.88 |microJy             |3.81E+13|  1.46E-05|+/-8.80E-07|Jy|2011AJ....141....1T|rms uncertainty|     7.872 microns   | Broad-band measurement|189.367981 62.315258 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
6|16 microns (IRS)    | 55.0      |+/-9.4  |microJy             |1.90E+13|  5.50E-05|+/-9.40E-06|Jy|2011AJ....141....1T|rms uncertainty|      15.8 microns   | Broad-band measurement|189.367981 62.315258 (J2000)| From fitting to map|                                        |From new raw data
7|24 microns (MIPS)   | 48.4      |+/-5.2  |microJy             |1.27E+13|  4.84E-05|+/-5.20E-06|Jy|2011AJ....141....1T|rms uncertainty|     23.68 microns   | Broad-band measurement|189.367981 62.315258 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
8|24 microns (MIPS)   | 54.8      |+/-3.1  |microJy             |1.27E+13|  5.48E-05|+/-3.10E-06|Jy|2011A&A...528A..35M|uncertainty|     23.68 microns   | Broad-band measurement|12 37 28.32 +62 18 54.86 (J2000)| Flux integrated from map|                                        |From new raw data
9|70 microns (MIPS)   ||<4.6       |milliJy             |4.20E+12||4.60E-03|Jy|2011A&A...528A..35M|no uncertainty reported|     71.42 microns   | Broad-band measurement|12 37 28.32 +62 18 54.86 (J2000)| Flux integrated from map|                                        |From new raw data
8|1.4 GHz (VLA)       | 37.2      |+/-11.1 |microJy             |1.40E+09|  3.72E-05|+/-1.11E-05|Jy|2010ApJS..188..178M|uncertainty|       1.4 GHz       | Broad-band measurement|12 37 28.34 +62 18 55.1 (J2000)| Total flux; Beam filling or dilution corrected|Major=2.1"; Minor=0.2"; PA=173 deg      |From new raw data
9|1.4 GHz (VLA)       | 46        |+/-8    | microJy            |1.40E+09|  4.60E-05|+/-8.00E-06|Jy|2006MNRAS.371..963B|1 sigma|       1.4 GHz       | Broad-band measurement|12 37 28.337 +62 18 54.79 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
10|1.4 GHz (VLA)       | 28        |+/-10    | microJy            |1.40E+09|  2.80E-05|+/-10.0E-06|Jy|2006MNRAS.371..963B|1 sigma|       1.4 GHz       | Broad-band measurement|12 37 28.337 +62 18 54.79 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
12|1.4 GHz (VLA)       | 37.2      |+/-11.1 |microJy             |1.40E+09|  3.72E-05|+/-1.11E-05|Jy|2010ApJS..188..178M|uncertainty|       1.4 GHz       | Broad-band measurement|12 37 28.34 +62 18 55.1 (J2000)| Total flux; Beam filling or dilution corrected|Major=2.1"; Minor=0.2"; PA=173 deg      |From new raw data
