
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2017-01-03T03:36:10PST



Photometric Data for SDSS J102434.56+470909.5

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|2-5 keV (XMM)       | 0.9E-15   ||erg/cm^2^/s         |8.46E+17|  1.06E-10||Jy|2010NewA...15...58I|no uncertainty reported|      3.50 keV       | Broad-band measurement|10 24 34.57 +47 09 09.9 (J2000)| Modelled datum|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
2|0.5-2 keV (XMM)     | 1.3E-15   ||erg/cm^2^/s         |3.02E+17|  4.30E-10||Jy|2010NewA...15...58I|no uncertainty reported|      1.25 keV       | Broad-band measurement|10 24 34.57 +47 09 09.9 (J2000)| Modelled datum|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
3|u (SDSS PSF) AB     | 21.710    |+/-0.214|asinh mag           |8.36E+14|  7.76E-06|+/-1.54E-06|Jy|2007SDSS6.C...0000:|based on count statistics only|3585       A         | Broad-band measurement|156.1440032823 47.1526651398 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; ELLIPFAINT - no isophotal fits performed; BINNED1 - detected at >=5 sigma in original imaging frame;|From new raw data
4|u (SDSS CModel) AB  | 21.815    ||asinh mag           |8.36E+14|  7.04E-06||Jy|2007SDSS6.C...0000:|no uncertainty reported|3585       A         | Broad-band measurement|156.1440032823 47.1526651398 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; ELLIPFAINT - no isophotal fits performed; BINNED1 - detected at >=5 sigma in original imaging frame;|From new raw data
5|u (SDSS Model) AB   | 21.801    |+/-0.248|asinh mag           |8.36E+14|  7.13E-06|+/-1.65E-06|Jy|2007SDSS6.C...0000:|based on count statistics only|3585       A         | Broad-band measurement|156.1440032823 47.1526651398 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; ELLIPFAINT - no isophotal fits performed; BINNED1 - detected at >=5 sigma in original imaging frame;|From new raw data
6|g (SDSS PSF) AB     | 21.298    |+/-0.055|asinh mag           |6.17E+14|  1.10E-05|+/-5.57E-07|Jy|2007SDSS6.C...0000:|based on count statistics only|4858       A         | Broad-band measurement|156.1440032823 47.1526651398 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
7|g (SDSS CModel) AB  | 21.202    ||asinh mag           |6.17E+14|  1.20E-05||Jy|2007SDSS6.C...0000:|no uncertainty reported|4858       A         | Broad-band measurement|156.1440032823 47.1526651398 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
8|g (SDSS Model) AB   | 21.251    |+/-0.049|asinh mag           |6.17E+14|  1.15E-05|+/-5.18E-07|Jy|2007SDSS6.C...0000:|based on count statistics only|4858       A         | Broad-band measurement|156.1440032823 47.1526651398 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
9|r (SDSS CModel) AB  | 20.936    ||asinh mag           |4.77E+14|  1.53E-05||Jy|2007SDSS6.C...0000:|no uncertainty reported|6290       A         | Broad-band measurement|156.1440032823 47.1526651398 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding; CANONICAL_BAND - this band was primary (usually r);|From new raw data
10|r (SDSS PSF) AB     | 20.996    |+/-0.045|asinh mag           |4.77E+14|  1.45E-05|+/-6.02E-07|Jy|2007SDSS6.C...0000:|based on count statistics only|6290       A         | Broad-band measurement|156.1440032823 47.1526651398 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding; CANONICAL_BAND - this band was primary (usually r);|From new raw data
11|r (SDSS Model) AB   | 20.935    |+/-0.046|asinh mag           |4.77E+14|  1.53E-05|+/-6.51E-07|Jy|2007SDSS6.C...0000:|based on count statistics only|6290       A         | Broad-band measurement|156.1440032823 47.1526651398 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding; CANONICAL_BAND - this band was primary (usually r);|From new raw data
12|i (SDSS PSF) AB     | 20.570    |+/-0.050|asinh mag           |3.89E+14|  2.15E-05|+/-9.90E-07|Jy|2007SDSS6.C...0000:|based on count statistics only|7706       A         | Broad-band measurement|156.1440032823 47.1526651398 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
13|i (SDSS CModel) AB  | 20.052    ||asinh mag           |3.89E+14|  3.46E-05||Jy|2007SDSS6.C...0000:|no uncertainty reported|7706       A         | Broad-band measurement|156.1440032823 47.1526651398 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
14|i (SDSS Model) AB   | 20.477    |+/-0.049|asinh mag           |3.89E+14|  2.34E-05|+/-1.06E-06|Jy|2007SDSS6.C...0000:|based on count statistics only|7706       A         | Broad-band measurement|156.1440032823 47.1526651398 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
15|z (SDSS CModel) AB  | 19.734    ||asinh mag           |3.25E+14|  4.54E-05||Jy|2007SDSS6.C...0000:|no uncertainty reported|9222       A         | Broad-band measurement|156.1440032823 47.1526651398 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
16|z (SDSS PSF) AB     | 20.302    |+/-0.117|asinh mag           |3.25E+14|  2.67E-05|+/-2.94E-06|Jy|2007SDSS6.C...0000:|based on count statistics only|9222       A         | Broad-band measurement|156.1440032823 47.1526651398 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
17|z (SDSS Model) AB   | 20.203    |+/-0.119|asinh mag           |3.25E+14|  2.93E-05|+/-3.27E-06|Jy|2007SDSS6.C...0000:|based on count statistics only|9222       A         | Broad-band measurement|156.1440032823 47.1526651398 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
18|J (2MASS)           | 18.650    |+/-0.150| mag                |2.40E+14|  5.52E-05|+/-7.63E-06|Jy|2009MNRAS.393.1408C|uncertainty|      1.25 microns   | Broad-band measurement|10 24 34.50 +47 09 11.0 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
19|H (2MASS)           | 17.150    |+/-0.100| mag                |1.82E+14|  1.41E-04|+/-1.30E-05|Jy|2009MNRAS.393.1408C|uncertainty|      1.65 microns   | Broad-band measurement|10 24 34.50 +47 09 11.0 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
20|K (2MASS)           | 16.370    |+/-0.100| mag                |1.38E+14|  1.89E-04|+/-1.74E-05|Jy|2009MNRAS.393.1408C|uncertainty|      2.17 microns   | Broad-band measurement|10 24 34.50 +47 09 11.0 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
21|3.6 microns (IRAC)  | 2.6274E+02|+/-1.9176E+00|microJy             |8.44E+13|  2.63E-04|+/-1.92E-06|Jy|2013SSTSLC4.2....0C|uncertainty|3.55       microns   | Broad-band measurement|| Flux in fixed aperture|3.8" aperture                           |From new raw data
22|3.6 microns (IRAC)  | 3.2271E+02|+/-2.5108E+00|microJy             |8.44E+13|  3.23E-04|+/-2.51E-06|Jy|2013SSTSLC4.2....0C|uncertainty|3.55       microns   | Broad-band measurement|| Flux in fixed aperture|5.8" aperture                           |From new raw data
23|4.5 microns (IRAC)  | 2.9126E+02|+/-2.7585E+00|microJy             |6.67E+13|  2.91E-04|+/-2.76E-06|Jy|2013SSTSLC4.2....0C|uncertainty|4.493      microns   | Broad-band measurement|| Flux in fixed aperture|3.8" aperture                           |From new raw data
24|4.5 microns (IRAC)  | 3.4244E+02|+/-3.3433E+00|microJy             |6.67E+13|  3.42E-04|+/-3.34E-06|Jy|2013SSTSLC4.2....0C|uncertainty|4.493      microns   | Broad-band measurement|| Flux in fixed aperture|5.8" aperture                           |From new raw data
25|5.8 microns (IRAC)  | 4.0658E+02|+/-1.4643E+01|microJy             |5.23E+13|  4.07E-04|+/-1.46E-05|Jy|2013SSTSLC4.2....0C|uncertainty|5.731      microns   | Broad-band measurement|| Flux in fixed aperture|5.8" aperture                           |From new raw data
26|5.8 microns (IRAC)  | 4.2040E+02|+/-1.0979E+01|microJy             |5.23E+13|  4.20E-04|+/-1.10E-05|Jy|2013SSTSLC4.2....0C|uncertainty|5.731      microns   | Broad-band measurement|| Flux in fixed aperture|3.8" aperture                           |From new raw data
27|8.0 microns (IRAC)  | 9.2297E+02|+/-1.2093E+01|microJy             |3.81E+13|  9.23E-04|+/-1.21E-05|Jy|2013SSTSLC4.2....0C|uncertainty|7.872      microns   | Broad-band measurement|| Flux in fixed aperture|5.8" aperture                           |From new raw data
28|8.0 microns (IRAC)  | 9.1978E+02|+/-9.6903E+00|microJy             |3.81E+13|  9.20E-04|+/-9.69E-06|Jy|2013SSTSLC4.2....0C|uncertainty|7.872      microns   | Broad-band measurement|| Flux in fixed aperture|3.8" aperture                           |From new raw data
29|12 microns (IRAS)   ||<8.305E-02 |Jy                  |2.50E+13||8.31E-02|Jy|1990IRASF.C...0000M|90% confidence| 12        microns   | Broad-band measurement|102129.9 +472442 (B1950)| Flux in fixed aperture|                                        |From new raw data
30|25 microns (IRAS)   ||<1.279E-01 |Jy                  |1.20E+13||1.28E-01|Jy|1990IRASF.C...0000M|90% confidence| 25        microns   | Broad-band measurement|102129.9 +472442 (B1950)| Flux in fixed aperture|                                        |From new raw data
31|[O IV] (Herschel)   ||<6E-18     |W/m^2^              |1.15E+13||6.00E+08|Jy-Hz|2010A&A...518L..36S|no uncertainty reported|        26 microns   | Line measurement; flux integrated over line; lines measured in emission|| From fitting to map|                                        |From new raw data
32|[S III] (Herschel)  ||<3E-18     |W/m^2^              |9.08E+12||3.00E+08|Jy-Hz|2010A&A...518L..36S|no uncertainty reported|        33 microns   | Line measurement; flux integrated over line; lines measured in emission|| From fitting to map|                                        |From new raw data
33|[O III] (Herschel)  | 0.9E-18   |+/-0.3E-18|W/m^2^              |5.77E+12|  9.00E+07|+/-3.00E+07|Jy-Hz|2010A&A...518L..36S|uncertainty|        52 microns   | Line measurement; flux integrated over line; lines measured in emission|| From fitting to map|                                        |From new raw data
34|60 microns (IRAS)   | 2.046E-01 |+/-22  %|Jy                  |5.00E+12|  2.05E-01|+/-4.50E-02|Jy|1990IRASF.C...0000M|uncertainty| 60        microns   | Broad-band measurement|102129.9 +472442 (B1950)| Flux in fixed aperture|IRAS quality flag = 3                   |From new raw data
35|100 microns (IRAS)  | 5.733E-01 |+/-24  %|Jy                  |3.00E+12|  5.73E-01|+/-1.38E-01|Jy|1990IRASF.C...0000M|uncertainty| 100       microns   | Broad-band measurement|102129.9 +472442 (B1950)| Flux in fixed aperture|IRAS quality flag = 2                   |From new raw data
36|350 microns (SHARC) | 0.383     |+/-0.051|Jy                  |8.57E+11|  3.83E-01|+/-5.10E-02|Jy|1999CIT...T00R....B|1 sigma|350        microns   | Broad-band measurement|102131.1 +472423. (B1950)| Flux integrated from map|                                        |From new raw data; OBJ_NAME modified from published value
37|CO(1-0) (GBT)       | 0.337     |+/-0.045|Jy km/s             |1.15E+11|  3.94E+04|+/-5.27E+03|Jy-Hz|2011ApJ...739L..32R|uncertainty|   115.271 GHz       | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|Measured with Spectrometer backend      |From new raw data
38|CO(1-0) (EVLA)      | 0.434     |+/-0.047|Jy km/s             |1.15E+11|  5.08E+04|+/-5.50E+03|Jy-Hz|2011ApJ...739L..32R|uncertainty|   115.271 GHz       | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|                                        |From new raw data
39|HCN(1-0) (GBT)      | 0.05      |+/-0.01 | Jy km/s            |8.86E+10|  4.50E+03|+/-9.00E+02|Jy-Hz|2004ApJ...614L..97V|uncertainty|     88.63 GHz       | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|S/N=5sigma                              |From new raw data
