
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-06-16T05:49:47PDT



Photometric Data for SDSS J141855.79+524749.3

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|u (SDSS PSF) AB     | 23.530    |+/-0.827|asinh mag           |8.36E+14|  1.27E-06|+/-1.26E-06|Jy|2007SDSS6.C...0000:|based on count statistics only|3585       A         | Broad-band measurement|214.7324700153 52.7970537858 (J2000)| Modelled datum|SDSS flags: CANONICAL_CENTER - used canonical, not local, center; NOPETRO - no Petrosian radius could be determined; NOPETRO_BIG - Petrosian radius is larger than extracted radial profile; BAD_RADIAL - some low S/N radial points; INTERP - object contains interpolated-over pixels; ELLIPFAINT - no isophotal fits performed; PSF_FLUX_INTERP - a signifcant amount of PSF's flux is interpolated; AMOMENT_FAINT - too faint for adaptive moments;|From new raw data
2|u (SDSS CModel) AB  | 21.720    ||asinh mag           |8.36E+14|  7.69E-06||Jy|2007SDSS6.C...0000:|no uncertainty reported|3585       A         | Broad-band measurement|214.7324700153 52.7970537858 (J2000)| Modelled datum|SDSS flags: CANONICAL_CENTER - used canonical, not local, center; NOPETRO - no Petrosian radius could be determined; NOPETRO_BIG - Petrosian radius is larger than extracted radial profile; BAD_RADIAL - some low S/N radial points; INTERP - object contains interpolated-over pixels; ELLIPFAINT - no isophotal fits performed; PSF_FLUX_INTERP - a signifcant amount of PSF's flux is interpolated; AMOMENT_FAINT - too faint for adaptive moments;|From new raw data
3|u (SDSS Model) AB   | 22.895    |+/-0.978|asinh mag           |8.36E+14|  2.51E-06|+/-2.45E-06|Jy|2007SDSS6.C...0000:|based on count statistics only|3585       A         | Broad-band measurement|214.7324700153 52.7970537858 (J2000)| Modelled datum|SDSS flags: CANONICAL_CENTER - used canonical, not local, center; NOPETRO - no Petrosian radius could be determined; NOPETRO_BIG - Petrosian radius is larger than extracted radial profile; BAD_RADIAL - some low S/N radial points; INTERP - object contains interpolated-over pixels; ELLIPFAINT - no isophotal fits performed; PSF_FLUX_INTERP - a signifcant amount of PSF's flux is interpolated; AMOMENT_FAINT - too faint for adaptive moments;|From new raw data
4|g (SDSS PSF) AB     | 23.939    |+/-0.421|asinh mag           |6.17E+14|  8.54E-07|+/-4.17E-07|Jy|2007SDSS6.C...0000:|based on count statistics only|4858       A         | Broad-band measurement|214.7324700153 52.7970537858 (J2000)| Modelled datum|SDSS flags: CANONICAL_CENTER - used canonical, not local, center; NOPETRO - no Petrosian radius could be determined; BAD_RADIAL - some low S/N radial points; PETROFAINT - Petrosian radius measured at very low surface brightness; ELLIPFAINT - no isophotal fits performed; AMOMENT_FAINT - too faint for adaptive moments;|From new raw data
5|g (SDSS CModel) AB  | 23.884    ||asinh mag           |6.17E+14|  9.10E-07||Jy|2007SDSS6.C...0000:|no uncertainty reported|4858       A         | Broad-band measurement|214.7324700153 52.7970537858 (J2000)| Modelled datum|SDSS flags: CANONICAL_CENTER - used canonical, not local, center; NOPETRO - no Petrosian radius could be determined; BAD_RADIAL - some low S/N radial points; PETROFAINT - Petrosian radius measured at very low surface brightness; ELLIPFAINT - no isophotal fits performed; AMOMENT_FAINT - too faint for adaptive moments;|From new raw data
6|g (SDSS Model) AB   | 23.329    |+/-0.758|asinh mag           |6.17E+14|  1.63E-06|+/-1.23E-06|Jy|2007SDSS6.C...0000:|based on count statistics only|4858       A         | Broad-band measurement|214.7324700153 52.7970537858 (J2000)| Modelled datum|SDSS flags: CANONICAL_CENTER - used canonical, not local, center; NOPETRO - no Petrosian radius could be determined; BAD_RADIAL - some low S/N radial points; PETROFAINT - Petrosian radius measured at very low surface brightness; ELLIPFAINT - no isophotal fits performed; AMOMENT_FAINT - too faint for adaptive moments;|From new raw data
7|r (SDSS CModel) AB  | 21.401    ||asinh mag           |4.77E+14|  9.97E-06||Jy|2007SDSS6.C...0000:|no uncertainty reported|6290       A         | Broad-band measurement|214.7324700153 52.7970537858 (J2000)| Modelled datum|SDSS flags: NOPETRO - no Petrosian radius could be determined; BAD_RADIAL - some low S/N radial points; PETROFAINT - Petrosian radius measured at very low surface brightness; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding; CANONICAL_BAND - this band was primary (usually r); AMOMENT_FAINT - too faint for adaptive moments; AMOMENT_MAXITER - too many iterations while determining adaptive moments;|From new raw data
8|r (SDSS PSF) AB     | 22.632    |+/-0.166|asinh mag           |4.77E+14|  3.16E-06|+/-5.01E-07|Jy|2007SDSS6.C...0000:|based on count statistics only|6290       A         | Broad-band measurement|214.7324700153 52.7970537858 (J2000)| Modelled datum|SDSS flags: NOPETRO - no Petrosian radius could be determined; BAD_RADIAL - some low S/N radial points; PETROFAINT - Petrosian radius measured at very low surface brightness; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding; CANONICAL_BAND - this band was primary (usually r); AMOMENT_FAINT - too faint for adaptive moments; AMOMENT_MAXITER - too many iterations while determining adaptive moments;|From new raw data
9|r (SDSS Model) AB   | 21.401    |+/-0.166|asinh mag           |4.77E+14|  9.97E-06|+/-1.53E-06|Jy|2007SDSS6.C...0000:|based on count statistics only|6290       A         | Broad-band measurement|214.7324700153 52.7970537858 (J2000)| Modelled datum|SDSS flags: NOPETRO - no Petrosian radius could be determined; BAD_RADIAL - some low S/N radial points; PETROFAINT - Petrosian radius measured at very low surface brightness; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding; CANONICAL_BAND - this band was primary (usually r); AMOMENT_FAINT - too faint for adaptive moments; AMOMENT_MAXITER - too many iterations while determining adaptive moments;|From new raw data
10|i (SDSS PSF) AB     | 22.976    |+/-0.319|asinh mag           |3.89E+14|  2.16E-06|+/-7.42E-07|Jy|2007SDSS6.C...0000:|based on count statistics only|7706       A         | Broad-band measurement|214.7324700153 52.7970537858 (J2000)| Modelled datum|SDSS flags: CANONICAL_CENTER - used canonical, not local, center; BAD_RADIAL - some low S/N radial points; ELLIPFAINT - no isophotal fits performed; AMOMENT_FAINT - too faint for adaptive moments;|From new raw data
11|i (SDSS CModel) AB  | 21.810    ||asinh mag           |3.89E+14|  6.79E-06||Jy|2007SDSS6.C...0000:|no uncertainty reported|7706       A         | Broad-band measurement|214.7324700153 52.7970537858 (J2000)| Modelled datum|SDSS flags: CANONICAL_CENTER - used canonical, not local, center; BAD_RADIAL - some low S/N radial points; ELLIPFAINT - no isophotal fits performed; AMOMENT_FAINT - too faint for adaptive moments;|From new raw data
12|i (SDSS Model) AB   | 21.513    |+/-0.283|asinh mag           |3.89E+14|  8.96E-06|+/-2.36E-06|Jy|2007SDSS6.C...0000:|based on count statistics only|7706       A         | Broad-band measurement|214.7324700153 52.7970537858 (J2000)| Modelled datum|SDSS flags: CANONICAL_CENTER - used canonical, not local, center; BAD_RADIAL - some low S/N radial points; ELLIPFAINT - no isophotal fits performed; AMOMENT_FAINT - too faint for adaptive moments;|From new raw data
13|z (SDSS PSF) AB     | 21.285    |+/-0.259|asinh mag           |3.25E+14|  1.03E-05|+/-2.76E-06|Jy|2007SDSS6.C...0000:|based on count statistics only|9222       A         | Broad-band measurement|214.7324700153 52.7970537858 (J2000)| Modelled datum|SDSS flags: CANONICAL_CENTER - used canonical, not local, center; BAD_RADIAL - some low S/N radial points; PETROFAINT - Petrosian radius measured at very low surface brightness; ELLIPFAINT - no isophotal fits performed; AMOMENT_FAINT - too faint for adaptive moments;|From new raw data
14|z (SDSS CModel) AB  | 20.668    ||asinh mag           |3.25E+14|  1.89E-05||Jy|2007SDSS6.C...0000:|no uncertainty reported|9222       A         | Broad-band measurement|214.7324700153 52.7970537858 (J2000)| Modelled datum|SDSS flags: CANONICAL_CENTER - used canonical, not local, center; BAD_RADIAL - some low S/N radial points; PETROFAINT - Petrosian radius measured at very low surface brightness; ELLIPFAINT - no isophotal fits performed; AMOMENT_FAINT - too faint for adaptive moments;|From new raw data
15|z (SDSS Model) AB   | 20.124    |+/-0.275|asinh mag           |3.25E+14|  3.16E-05|+/-8.11E-06|Jy|2007SDSS6.C...0000:|based on count statistics only|9222       A         | Broad-band measurement|214.7324700153 52.7970537858 (J2000)| Modelled datum|SDSS flags: CANONICAL_CENTER - used canonical, not local, center; BAD_RADIAL - some low S/N radial points; PETROFAINT - Petrosian radius measured at very low surface brightness; ELLIPFAINT - no isophotal fits performed; AMOMENT_FAINT - too faint for adaptive moments;|From new raw data
16|K_s (Keck)          | 17.59     || mag                |1.39E+14|  5.71E-05||Jy|2007MNRAS.382..109T|no uncertainty reported|      2.15 microns   | Broad-band measurement|214.73238 +52.79687 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
