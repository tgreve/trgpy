
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-07-08T06:57:45PDT



Photometric Data for GOODS J123718.58+621315.4

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|U (KPNO) AB         | 24.11     ||mag                 |8.44E+14|  8.24E-07||Jy|2006ApJ...653.1004R|no uncertainty reported|    3550   A         | Broad-band measurement|123718.58 +621315.0 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data; derived from aflux in a different band and a color
2|U (KPNO) AB         | 23.9      || mag                |8.22E+14|  1.00E-06||Jy|2004AJ....127.3137C|no uncertainty reported| 3647.65   A         | Broad-band measurement|189.327408 +62.22095 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
3|B F435W (HST/ACS) AB      | 23.585    ||mag                 |6.98E+14|  1.34E-06||Jy|2007ApJ...660...81M|no uncertainty reported|    4297   A         | Broad-band measurement|12 37 18.564 +62 13 15.06 (J2000)| Flux integrated from map|                                        |From reprocessed raw data; Corrected for contaminatingsources
4|B (Subaru) AB       | 23.64     ||mag                 |6.77E+14|  1.27E-06||Jy|2006ApJ...653.1027W|no uncertainty reported| 4427.60   A         | Broad-band measurement|189.327350 62.220850 (J2000)| Flux in fixed aperture|3" diameter aperture                    |Averaged from previously published data
5|B (Subaru) AB       | 23.6      || mag                |6.77E+14|  1.32E-06||Jy|2004AJ....127.3137C|no uncertainty reported| 4427.60   A         | Broad-band measurement|189.327408 +62.22095 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
6|G (KECK) AB         | 23.63     ||mag                 |6.27E+14|  1.28E-06||Jy|2006ApJ...653.1004R|no uncertainty reported|    4780   A         | Broad-band measurement|123718.58 +621315.0 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data; derived from aflux in a different band and a color
7|V (Subaru) AB       | 23.6      || mag                |5.48E+14|  1.32E-06||Jy|2004AJ....127.3137C|no uncertainty reported| 5471.22   A         | Broad-band measurement|189.327408 +62.22095 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
8|V (HST/ACS) AB      | 23.360    ||mag                 |5.08E+14|  1.64E-06||Jy|2007ApJ...660...81M|no uncertainty reported|    5907   A         | Broad-band measurement|12 37 18.564 +62 13 15.06 (J2000)| Flux integrated from map|                                        |From reprocessed raw data; Corrected for contaminatingsources
9|R (Keck II) AB      | 23.54     || mag                |4.62E+14|  1.39E-06||Jy|2004AJ....127.3121W|no uncertainty reported|   648.7   A         | Broad-band measurement|12 37 18.564 +62 13 15.06 (J2000)| Total flux|                                        |From new raw data
10|R (Subaru) AB       | 23.37     ||mag                 |4.59E+14|  1.63E-06||Jy|2006ApJ...653.1027W|no uncertainty reported| 6534.16   A         | Broad-band measurement|189.327350 62.220850 (J2000)| Flux in fixed aperture|3" diameter aperture                    |Averaged from previously published data
11|R (Subaru) AB       | 23.4      || mag                |4.59E+14|  1.59E-06||Jy|2004AJ....127.3137C|no uncertainty reported| 6534.16   A         | Broad-band measurement|189.327408 +62.22095 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
12|R (KECK) AB         | 23.35     ||mag                 |4.39E+14|  1.66E-06||Jy|2006ApJ...653.1004R|no uncertainty reported|    6830   A         | Broad-band measurement|123718.58 +621315.0 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data
13|i F775W (HST/ACS) AB      | 23.089    ||mag                 |3.86E+14|  2.11E-06||Jy|2007ApJ...660...81M|no uncertainty reported|    7764   A         | Broad-band measurement|12 37 18.564 +62 13 15.06 (J2000)| Flux integrated from map|                                        |From reprocessed raw data; Corrected for contaminatingsources
14|I (Subaru) AB       | 23.17     ||mag                 |3.76E+14|  1.96E-06||Jy|2006ApJ...653.1027W|no uncertainty reported| 7975.89   A         | Broad-band measurement|189.327350 62.220850 (J2000)| Flux in fixed aperture|3" diameter aperture                    |Averaged from previously published data
15|I (Subaru) AB       | 23.2      || mag                |3.76E+14|  1.91E-06||Jy|2004AJ....127.3137C|no uncertainty reported| 7975.89   A         | Broad-band measurement|189.327408 +62.22095 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
16|z' (Subaru) AB      | 22.9      || mag                |3.31E+14|  2.51E-06||Jy|2004AJ....127.3137C|no uncertainty reported| 9069.21   A         | Broad-band measurement|189.327408 +62.22095 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
17|z F850LP (HST/ACS) AB      | 22.791    ||mag                 |3.17E+14|  2.78E-06||Jy|2007ApJ...660...81M|no uncertainty reported|    9445   A         | Broad-band measurement|12 37 18.564 +62 13 15.06 (J2000)| Flux integrated from map|                                        |From reprocessed raw data; Corrected for contaminatingsources
18|J (WIRC) AB         | 22.19     ||mag                 |2.40E+14|  4.83E-06||Jy|2006ApJ...653.1004R|no uncertainty reported|   1.250   microns   | Broad-band measurement|123718.58 +621315.0 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data
19|HK' (UH) AB         | 22.2      || mag                |1.58E+14|  4.79E-06||Jy|2004AJ....127.3137C|no uncertainty reported|18947.38   A         | Broad-band measurement|189.327408 +62.22095 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
20|HK' (QUIRC) AB      | 22.19     |+/-0.29 |mag                 |1.58E+14|  4.83E-06|+/-1.29E-06|Jy|2006ApJ...653.1027W|uncertainty|18947.38   A         | Broad-band measurement|189.327350 62.220850 (J2000)| Flux in fixed aperture|3" diameter aperture                    |Averaged from previously published data
21|K_s (WIRC) AB       | 21.94     ||mag                 |1.39E+14|  6.08E-06||Jy|2006ApJ...653.1004R|no uncertainty reported|   2.150   microns   | Broad-band measurement|123718.58 +621315.0 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data
22|3.6 microns IRAC AB | 21.75     |+/-0.07 |mag                 |8.44E+13|  7.25E-06|+/-4.67E-07|Jy|2006ApJ...653.1004R|uncertainty|   3.550   microns   | Broad-band measurement|123718.58 +621315.0 (J2000)| Flux integrated from map|                                        |From new raw data
23|4.5 microns IRAC AB | 21.72     |+/-0.07 |mag                 |6.67E+13|  7.45E-06|+/-4.80E-07|Jy|2006ApJ...653.1004R|uncertainty|   4.493   microns   | Broad-band measurement|123718.58 +621315.0 (J2000)| Flux integrated from map|                                        |From new raw data
24|5.8 microns IRAC AB | 21.96     |+/-0.25 |mag                 |5.23E+13|  5.97E-06|+/-1.38E-06|Jy|2006ApJ...653.1004R|uncertainty|   5.731   microns   | Broad-band measurement|123718.58 +621315.0 (J2000)| Flux integrated from map|                                        |From new raw data
25|8.0 microns IRAC AB | 21.67     |+/-0.07 |mag                 |3.81E+13|  7.80E-06|+/-5.03E-07|Jy|2006ApJ...653.1004R|uncertainty|   7.872   microns   | Broad-band measurement|123718.58 +621315.0 (J2000)| Flux integrated from map|                                        |From new raw data
26|24 microns (MIPS)   | 64.8      |+/-8.3  |microJy             |1.27E+13|  6.48E-05|+/-8.30E-06|Jy|2006ApJ...653.1004R|uncertainty|   23.68   microns   | Broad-band measurement|123718.58 +621315.0 (J2000)| Flux integrated from map|                                        |From new raw data
27|24 microns (MIPS)   | 47.0      |+/-4.3  |microJy             |1.27E+13|  4.70E-05|+/-4.30E-06|Jy|2011A&A...528A..35M|uncertainty|     23.68 microns   | Broad-band measurement|12 37 18.58 +62 13 15.03 (J2000)| Flux integrated from map|                                        |From new raw data
1|24 microns (MIPS)   | 73.       |+/-23.   |microJy             |1.27E+13|73.E-06|+/-23.0E-06|Jy|2009ApJ...694.1517D|3sigma uncertainty|     23.68 microns   | Broad-band measurement|12 37 11.89 +62 22 11.8 (J2000)| Flux integrated from map|                                        |From new raw data
28|70 microns (MIPS)   ||<4.4       |milliJy             |4.20E+12||4.40E-03|Jy|2011A&A...528A..35M|no uncertainty reported|     71.42 microns   | Broad-band measurement|12 37 18.58 +62 13 15.03 (J2000)| Flux integrated from map|                                        |From new raw data
2|70 microns (MIPS)   |           |<2.6  |mJy             |4.20E+12| |2.6E-03|Jy|2009ApJ...699.1610H|3 sigma|     71.42 microns   | Broad-band measurement|221804.42 +002154.4 (J2000)| Flux in fixed aperture|                                        |From new raw data
3|850 microns (SCUBA) |           |<5.7    |mJy             |3.53E+11|  |5.7E-03|Jy|2005MNRAS.358..149P|3sigma uncertainty|     850   microns   | Broad-band measurement|12 37 11.7 +62 22 12 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
4|1200 microns (MAMBO)|           |<0.9    |mJy             |2.50E+11|        |0.9E-03|Jy|2004MNRAS.354..779G|3rms uncertainty|      1200 microns   | Broad-band measurement|16 36 55.9 +40 59 12 (J2000)| Flux integrated from map|S/N = 3.66                              |From new raw data
5|1.4 GHz (VLA)       | 15.2     |+/-6.8  | microJy        |1.40E+09| 15.2E-06|+/-6.8E-06|Jy|2006MNRAS.371..963B|1 sigma|       1.4 GHz       | Broad-band measurement|16 36 55.767 +40 59 09.97 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
