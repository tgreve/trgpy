
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-07-08T02:08:52PDT



Photometric Data for ACS-GC 50012028

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
15|U (KPNO) AB         | 23.9      || mag                |8.22E+14|  1.00E-06||Jy|2004AJ....127.3137C|no uncertainty reported| 3647.65   A         | Broad-band measurement|189.140244 +62.16839 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
16|B F435W (HST/ACS) AB      | 23.602    ||mag                 |6.98E+14|  1.32E-06||Jy|2007ApJ...660...81M|no uncertainty reported|    4297   A         | Broad-band measurement|12 36 33.637 +62 10 05.89 (J2000)| Flux integrated from map|                                        |From reprocessed raw data; Corrected for contaminatingsources
17|F435W (HST/ACS) AB      | 21.336    |+/-0.008|mag                 |6.92E+14|  1.06E-05|+/-7.82E-08|Jy|2011ApJ...734..121S|uncertainty|      4333 A         | Broad-band measurement|189.140244 62.168388 (J2000)| Total flux|                                        |From reprocessed raw data
18|F435W (HST/ACS) AB      | 26.40     |+/-0.30 |mag                 |6.92E+14|  1.00E-07|+/-2.76E-08|Jy|2011ApJ...734..121S|uncertainty|      4333 A         | Broad-band measurement|189.140244 62.168388 (J2000)| Modelled datum|Central point source mag                |From reprocessed raw data
19|F435W (HST/ACS) AB      | 21.35     |+/-0.19 |mag                 |6.92E+14|  1.05E-05|+/-1.83E-06|Jy|2011ApJ...734..121S|uncertainty|      4333 A         | Broad-band measurement|189.140244 62.168388 (J2000)| Modelled datum|Host galaxy mag                         |From reprocessed raw data
20|B (Subaru) AB       | 23.9      || mag                |6.77E+14|  1.00E-06||Jy|2004AJ....127.3137C|no uncertainty reported| 4427.60   A         | Broad-band measurement|189.140244 +62.16839 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
21|B (Subaru) AB       | 23.92     ||mag                 |6.77E+14|  9.82E-07||Jy|2006ApJ...653.1027W|no uncertainty reported| 4427.60   A         | Broad-band measurement|189.140154 62.168303 (J2000)| Flux in fixed aperture|3" diameter aperture                    |Averaged from previously published data
22|V (Subaru) AB       | 23.4      || mag                |5.48E+14|  1.59E-06||Jy|2004AJ....127.3137C|no uncertainty reported| 5471.22   A         | Broad-band measurement|189.140244 +62.16839 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
23|V (HST/ACS) AB      | 22.834    ||mag                 |5.08E+14|  2.67E-06||Jy|2007ApJ...660...81M|no uncertainty reported|    5907   A         | Broad-band measurement|12 36 33.637 +62 10 05.89 (J2000)| Flux integrated from map|                                        |From reprocessed raw data; Corrected for contaminatingsources
24|R (Keck II) AB      | 22.96     || mag                |4.62E+14|  2.38E-06||Jy|2004AJ....127.3121W|no uncertainty reported|   648.7   A         | Broad-band measurement|12 36 33.637 +62 10 05.89 (J2000)| Total flux|                                        |From new raw data
25|R (Subaru) AB       | 22.9      || mag                |4.59E+14|  2.51E-06||Jy|2004AJ....127.3137C|no uncertainty reported| 6534.16   A         | Broad-band measurement|189.140244 +62.16839 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
26|R (Subaru) AB       | 22.84     ||mag                 |4.59E+14|  2.65E-06||Jy|2006ApJ...653.1027W|no uncertainty reported| 6534.16   A         | Broad-band measurement|189.140154 62.168303 (J2000)| Flux in fixed aperture|3" diameter aperture                    |Averaged from previously published data
27|R (Subaru) AB       | 22.60     ||mag                 |4.58E+14|  3.31E-06||Jy|2007MNRAS.377..203G|no uncertainty reported|    6550   A         | Broad-band measurement|12 36 33.67 +62 10 05.7 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
28|i F775W (HST/ACS) AB      | 21.838    ||mag                 |3.86E+14|  6.68E-06||Jy|2007ApJ...660...81M|no uncertainty reported|    7764   A         | Broad-band measurement|12 36 33.637 +62 10 05.89 (J2000)| Flux integrated from map|                                        |From reprocessed raw data; Corrected for contaminatingsources
29|I (Subaru) AB       | 22.0      || mag                |3.76E+14|  5.75E-06||Jy|2004AJ....127.3137C|no uncertainty reported| 7975.89   A         | Broad-band measurement|189.140244 +62.16839 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
30|I (Subaru) AB       | 22.02     ||mag                 |3.76E+14|  5.65E-06||Jy|2006ApJ...653.1027W|no uncertainty reported| 7975.89   A         | Broad-band measurement|189.140154 62.168303 (J2000)| Flux in fixed aperture|3" diameter aperture                    |Averaged from previously published data
31|z' (Subaru) AB      | 21.7      || mag                |3.31E+14|  7.59E-06||Jy|2004AJ....127.3137C|no uncertainty reported| 9069.21   A         | Broad-band measurement|189.140244 +62.16839 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
32|z F850LP (HST/ACS) AB      | 21.308    ||mag                 |3.17E+14|  1.09E-05||Jy|2007ApJ...660...81M|no uncertainty reported|    9445   A         | Broad-band measurement|12 36 33.637 +62 10 05.89 (J2000)| Flux integrated from map|                                        |From reprocessed raw data; Corrected for contaminatingsources
33|HK' (UH) AB         | 20.3      || mag                |1.58E+14|  2.75E-05||Jy|2004AJ....127.3137C|no uncertainty reported|18947.38   A         | Broad-band measurement|189.140244 +62.16839 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
34|HK' (QUIRC) AB      | 20.26     |+/-0.06 |mag                 |1.58E+14|  2.86E-05|+/-1.58E-06|Jy|2006ApJ...653.1027W|uncertainty|18947.38   A         | Broad-band measurement|189.140154 62.168303 (J2000)| Flux in fixed aperture|3" diameter aperture                    |Averaged from previously published data
35|3.6 microns (IRAC)  | 74.20     |+/-3.71 |microJy             |8.44E+13|  7.42E-05|+/-3.71E-06|Jy|2011AJ....141....1T|rms uncertainty|     3.550 microns   | Broad-band measurement|189.140320 62.168324 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
36|3.6 microns (IRAC)  | 72.48     |+/-0.07 |microJy             |8.44E+13|  7.25E-05|+/-7.00E-08|Jy|2007MNRAS.377..203G|uncertainty|   3.550   microns   | Broad-band measurement|12 36 33.67 +62 10 05.7 (J2000)| Corrected to total flux from single aperture measurement|                                        |From reprocessed raw data
37|4.5 microns (IRAC)  | 56.80     |+/-2.84 |microJy             |6.67E+13|  5.68E-05|+/-2.84E-06|Jy|2011AJ....141....1T|rms uncertainty|     4.493 microns   | Broad-band measurement|189.140320 62.168324 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
38|4.5 microns (IRAC)  | 56.94     |+/-0.09 |microJy             |6.67E+13|  5.69E-05|+/-9.00E-08|Jy|2007MNRAS.377..203G|uncertainty|   4.493   microns   | Broad-band measurement|12 36 33.67 +62 10 05.7 (J2000)| Corrected to total flux from single aperture measurement|                                        |From reprocessed raw data
39|5.8 microns (IRAC)  | 44.90     |+/-2.29 |microJy             |5.23E+13|  4.49E-05|+/-2.29E-06|Jy|2011AJ....141....1T|rms uncertainty|     5.731 microns   | Broad-band measurement|189.140320 62.168324 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
40|5.8 microns (IRAC)  | 45.76     |+/-0.48 |microJy             |5.23E+13|  4.58E-05|+/-4.80E-07|Jy|2007MNRAS.377..203G|uncertainty|   5.731   microns   | Broad-band measurement|12 36 33.67 +62 10 05.7 (J2000)| Corrected to total flux from single aperture measurement|                                        |From reprocessed raw data
41|8.0 microns (IRAC)  | 48.24     |+/-0.53 |microJy             |3.81E+13|  4.82E-05|+/-5.30E-07|Jy|2007MNRAS.377..203G|uncertainty|   7.872   microns   | Broad-band measurement|12 36 33.67 +62 10 05.7 (J2000)| Corrected to total flux from single aperture measurement|                                        |From reprocessed raw data
42|8.0 microns (IRAC)  | 49.50     |+/-2.53 |microJy             |3.81E+13|  4.95E-05|+/-2.53E-06|Jy|2011AJ....141....1T|rms uncertainty|     7.872 microns   | Broad-band measurement|189.140320 62.168324 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
43|11 microns (AKARI)  | 94.0      |+/-15   | microJy            |2.73E+13|  9.40E-05|+/-1.50E-05|Jy|2009MNRAS.394..375N|uncertainty|        11 microns   | Broad-band measurement|12 36 33.66 +62 10 06.20 (J2000)| Flux integrated from map|                                        |From new raw data
44|16 microns (IRS)    | 528.4     |+/-14.8 |microJy             |1.90E+13|  5.28E-04|+/-1.48E-05|Jy|2011AJ....141....1T|rms uncertainty|      15.8 microns   | Broad-band measurement|189.140320 62.168324 (J2000)| From fitting to map|                                        |From new raw data
45|16 microns (IRS)    | 438       |+/-25   | microJy            |1.87E+13|  4.38E-04|+/-2.50E-05|Jy|2009MNRAS.394..375N|uncertainty|        16 microns   | Broad-band measurement|12 36 33.66 +62 10 06.20 (J2000)| Flux integrated from map|                                        |Averaged from previously published data
46|18 microns (AKARI)  | 398       |+/-32   | microJy            |1.67E+13|  3.98E-04|+/-3.20E-05|Jy|2009MNRAS.394..375N|uncertainty|        18 microns   | Broad-band measurement|12 36 33.66 +62 10 06.20 (J2000)| Flux integrated from map|                                        |From new raw data
47|24 microns (MIPS)   | 581       |+/-9    |microJy             |1.27E+13|  5.81E-04|+/-9.00E-06|Jy|2011ApJ...726...93R|uncertainty|     23.68 microns   | Broad-band measurement|12 36 33.67 +62 10 05.8 (J2000)| Not reported in paper|                                        |Averaged from previously published data
48|24 microns (MIPS)   | 546.62    |+/-4.99 |microJy             |1.27E+13|  5.47E-04|+/-4.99E-06|Jy|2007MNRAS.377..203G|uncertainty|   23.68   microns   | Broad-band measurement|12 36 33.67 +62 10 05.7 (J2000)| Corrected to total flux from single aperture measurement|                                        |From reprocessed raw data
49|24 microns (MIPS)   | 576.8     |+/-4.9  |microJy             |1.27E+13|  5.77E-04|+/-4.90E-06|Jy|2011A&A...528A..35M|uncertainty|     23.68 microns   | Broad-band measurement|12 36 33.68 +62 10 05.90 (J2000)| Flux integrated from map|                                        |From new raw data
50|24 microns (MIPS)   | 581.0     |+/-9.0  |microJy             |1.27E+13|  5.81E-04|+/-9.00E-06|Jy|2011AJ....141....1T|rms uncertainty|     23.68 microns   | Broad-band measurement|189.140320 62.168324 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
1|24 microns (MIPS)   | 527.      |+/-7.0 |mJy            |1.27E+13|527.E-03|+/-7.E-03|Jy|2009ApJ...694.1517D|1rms uncertainty|     23.68 microns   | Broad-band measurement|12 37 11.89 +62 22 11.8 (J2000)| Flux integrated from map|                                        |From new raw data
51|70 microns (MIPS)   | 3.0       |+/-0.3  |milliJy             |4.20E+12|  3.00E-03|+/-3.00E-04|Jy|2011A&A...528A..35M|uncertainty|     71.42 microns   | Broad-band measurement|12 36 33.68 +62 10 05.90 (J2000)| Flux integrated from map|                                        |From new raw data
2| 70 microns (PACS)   | 2.7       |+/-0.6 |mJy            |4.283e+12|2.7E-03|+/-0.6E-03 |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
3|100 microns (PACS)  | 8.5       |+/-0.3 |mJy            |2.998e+12|8.5E-03|+/-0.3E-03|Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
3|160 microns (PACS)  | 16.3      |+/-1.0 |mJy            |1.874e+12|16.3E-03|+/-1.0E-03 |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
4|250 microns (SPIRE) | 20.2      |+/-2.5 |mJy            |1.199e+12|20.2E-03|+/-2.5e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
5|350 microns (SPIRE) | 13.0      |+/-3.0 |mJy            |8.565e+11|13.0E-03|+/-3.0e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
6|500 microns (SPIRE) |           |<12.0  |mJy            |5.996e+11| |12.0E-03|Jy |2.40e+01 |3sigma |bla |-9.90e+01 |-9.90e+01 | NaN|
7|1160 microns (Penner)|           |<1.6  |mJy            |2.58442e+08| |1.6E-03|Jy |2.40e+01 |3sigma |bla |-9.90e+01 |-9.90e+01 | NaN|
52|1.4 GHz (VLA)       | 46        ||microJy             |1.40E+09|  4.60E-05||Jy|2005MNRAS.358.1159M|no uncertainty reported|     1.4   GHz       | Broad-band measurement|12 36 33.7269 +62 10 05.962 (J2000)| Flux integrated from map|                                        |From new raw data
53|1.4 GHz (VLA)       | 58.5      |+/-9.1  |microJy             |1.40E+09|  5.85E-05|+/-9.10E-06|Jy|2010ApJS..188..178M|uncertainty|       1.4 GHz       | Broad-band measurement|12 36 33.67 +62 10 05.8 (J2000)| Total flux; Beam filling or dilution corrected|Major=1.2"; Minor=0.9"; PA=101 deg      |From new raw data
54|1.4 GHz (VLA)       | 52        |+/-11   | microJy            |1.40E+09|  5.20E-05|+/-1.10E-05|Jy|2006MNRAS.371..963B|1 sigma|       1.4 GHz       | Broad-band measurement|12 36 33.708 +62 10 05.90 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
55|1.4 GHz (VLA)       | 46.5      |+/-8.1  |microJy             |1.40E+09|  4.65E-05|+/-8.10E-06|Jy|2000ApJ...533..611R|1 sigma|1.4        GHz       | Broad-band measurement; broad-band flux derived by integration over spectrum; synthetic band|123633.739 +621006.16 (J2000)| Flux integrated from map; Pointing and beam filling|                                        |From new raw data; Corrected for contaminating sources
