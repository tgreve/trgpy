
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2017-01-03T06:58:11PST



Photometric Data for 2MASSi J1205231-074232

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|0.5-2 keV (Chandra) | 8.50E-15  ||ergs cm^-2^ s^-1^   |3.02E+17|  2.81E-09||Jy|2005AJ....129.2519V|no uncertainty reported|    1.25   keV       | Broad-band measurement|| Flux integrated from map|Corr. for quantum eff. decay at low E   |From new raw data; Extinction-corrected for Milky Way; NEDfrequency assigned to mid-point of band in keV
2|0.5-2 keV (Chandra) | 6E-15     ||erg cm^-2^ s^-1^    |3.02E+17|  1.99E-09||Jy|2006ApJ...645L..97I|no uncertainty reported|1.25       keV       | Broad-band measurement|12 05 23.12 -07 42 32.5 (J2000)| Flux integrated from map|                                        |From reprocessed raw data; NED frequency assigned tomid-point of band in keV
3|Ly{alpha} (Subaru)  | 2.7E-16   ||ergs/s/cm^2^        |2.46E+15|  2.70E+07||Jy-Hz|2004AJ....128.2704O|no uncertainty reported|      1216 A         | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|Total flux                              |From new raw data
4|Ly{alpha} (Subaru)  | 6.5E-17   ||ergs/s/cm^2^        |2.46E+15|  6.50E+06||Jy-Hz|2004AJ....128.2704O|no uncertainty reported|      1216 A         | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|Nuclear flux                            |From new raw data
5|3.6 microns (IRAC)  | 4.5049E+02|+/-3.4275E-01|microJy             |8.44E+13|  4.50E-04|+/-3.43E-07|Jy|2013SSTSLC4.2....0C|uncertainty|3.55       microns   | Broad-band measurement|| Flux in fixed aperture|3.8" aperture                           |From new raw data
6|3.6 microns (IRAC)  | 4.4927E+02|+/-3.2310E-01|microJy             |8.44E+13|  4.49E-04|+/-3.23E-07|Jy|2013SSTSLC4.2....0C|uncertainty|3.55       microns   | Broad-band measurement|| Flux in fixed aperture|5.8" aperture                           |From new raw data
7|3.6 microns (IRAC)  | 0.461     |+/-0.001|milliJy             |8.44E+13|  4.61E-04|+/-1.00E-06|Jy|2006ApJ...641L..85H|estimated error|   3.550   microns   | Broad-band measurement|| Corrected to total flux from single aperture measurement|Absolute calibration uncertainty is 3-5%|From new raw data
8|4.5 microns (IRAC)  | 3.6946E+02|+/-3.5854E-01|microJy             |6.67E+13|  3.69E-04|+/-3.59E-07|Jy|2013SSTSLC4.2....0C|uncertainty|4.493      microns   | Broad-band measurement|| Flux in fixed aperture|3.8" aperture                           |From new raw data
9|4.5 microns (IRAC)  | 3.7755E+02|+/-3.7323E-01|microJy             |6.67E+13|  3.78E-04|+/-3.73E-07|Jy|2013SSTSLC4.2....0C|uncertainty|4.493      microns   | Broad-band measurement|| Flux in fixed aperture|5.8" aperture                           |From new raw data
10|4.5 microns (IRAC)  | 0.375     |+/-0.001|milliJy             |6.67E+13|  3.75E-04|+/-1.00E-06|Jy|2006ApJ...641L..85H|estimated error|   4.493   microns   | Broad-band measurement|| Corrected to total flux from single aperture measurement|Absolute calibration uncertainty is 3-5%|From new raw data
11|5.8 microns (IRAC)  | 4.1163E+02|+/-9.6095E-01|microJy             |5.23E+13|  4.12E-04|+/-9.61E-07|Jy|2013SSTSLC4.2....0C|uncertainty|5.731      microns   | Broad-band measurement|| Flux in fixed aperture|5.8" aperture                           |From new raw data
12|5.8 microns (IRAC)  | 4.0502E+02|+/-8.5212E-01|microJy             |5.23E+13|  4.05E-04|+/-8.52E-07|Jy|2013SSTSLC4.2....0C|uncertainty|5.731      microns   | Broad-band measurement|| Flux in fixed aperture|3.8" aperture                           |From new raw data
13|5.8 microns (IRAC)  | 0.410     |+/-0.001|milliJy             |5.23E+13|  4.10E-04|+/-1.00E-06|Jy|2006ApJ...641L..85H|estimated error|   5.731   microns   | Broad-band measurement|| Corrected to total flux from single aperture measurement|Absolute calibration uncertainty is 3-5%|From new raw data
14|8.0 microns (IRAC)  | 0.657     |+/-0.002|milliJy             |3.81E+13|  6.57E-04|+/-2.00E-06|Jy|2006ApJ...641L..85H|estimated error|   7.872   microns   | Broad-band measurement|| Corrected to total flux from single aperture measurement|Absolute calibration uncertainty is 3-5%|From new raw data
15|8.0 microns (IRAC)  | 6.3122E+02|+/-1.5837E+00|microJy             |3.81E+13|  6.31E-04|+/-1.58E-06|Jy|2013SSTSLC4.2....0C|uncertainty|7.872      microns   | Broad-band measurement|| Flux in fixed aperture|5.8" aperture                           |From new raw data
16|8.0 microns (IRAC)  | 6.4882E+02|+/-1.2593E+00|microJy             |3.81E+13|  6.49E-04|+/-1.26E-06|Jy|2013SSTSLC4.2....0C|uncertainty|7.872      microns   | Broad-band measurement|| Flux in fixed aperture|3.8" aperture                           |From new raw data
17|24 microns (MIPS)   | 2.37      |+/-0.24 |milliJy             |1.27E+13|  2.37E-03|+/-2.40E-04|Jy|2006ApJ...641L..85H|estimated error|   23.68   microns   | Broad-band measurement|| Corrected to total flux from single aperture measurement|Absolute calibration uncertainty is 10% |From new raw data
18|24 microns (MIPS)   | 5.0497E+03|+/-5.4182E+01|microJy             |1.27E+13|  5.05E-03|+/-5.42E-05|Jy|2013SSTSLC4.2....0C|uncertainty|23.68      microns   | Broad-band measurement|| Modelled datum|PSF fit                                 |From new raw data
19|24 microns (MIPS)   | 5.1785E+03|+/-4.8452E+01|microJy             |1.27E+13|  5.18E-03|+/-4.85E-05|Jy|2013SSTSLC4.2....0C|uncertainty|23.68      microns   | Broad-band measurement|| Flux in fixed aperture|14.7" aperture                          |From new raw data
20|70 microns (PACS)   | 15.0      |+/-2.0  |milliJy             |4.28E+12|  1.50E-02|+/-2.00E-03|Jy|2010A&A...518L..34L|uncertainty|      70.0 microns   | Broad-band measurement|| Flux in fixed aperture|7.0" radius aperture                    |From new raw data
21|160 microns (PACS)  | 39.8      |+/-3.7  |milliJy             |1.87E+12|  3.98E-02|+/-3.70E-03|Jy|2010A&A...518L..34L|uncertainty|     160.0 microns   | Broad-band measurement|| Flux in fixed aperture|10.0" radius aperture                   |From new raw data
22|350 microns (SHARC-II)  | 0.106     |+/-0.007|Jy                  |8.57E+11|  1.06E-01|+/-7.00E-03|Jy|1999CIT...T00R....B|1 sigma|350        microns   | Broad-band measurement|120249.3 -072550. (B1950)| Flux integrated from map|                                        |From new raw data
23|870 microns (SMA)   | 32        |+/-4    |milliJy             |3.33E+11|  3.20E-02|+/-4.00E-03|Jy|2006ApJ...645L..97I|uncertainty| 900       microns   | Broad-band measurement|12 05 23.12 -07 42 32.5 (J2000)| Flux integrated from map|Beam size = 3.4" x 2.7"                 |From new raw data
24|1.25 mm (MAMBO)      | 10.5      |+/-1.5  |milliJy             |2.40E+11|  1.05E-02|+/-1.50E-03|Jy|1994MNRAS.267L...9M|estimated error|    1.25   mm        | Broad-band measurement|| Total flux|                                        |From new raw data
