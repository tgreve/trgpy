
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-07-08T05:26:23PDT



Photometric Data for ACS-GC 50000760

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|B F435W (HST/ACS) AB      | 22.968    ||mag                 |6.98E+14|  2.36E-06||Jy|2007ApJ...660...81M|no uncertainty reported|    4297   A         | Broad-band measurement|12 37 59.473 +62 17 33.06 (J2000)| Flux integrated from map|                                        |From reprocessed raw data; Corrected for contaminatingsources
2|B (Subaru) AB       | 23.47     ||mag                 |6.77E+14|  1.49E-06||Jy|2006ApJ...653.1027W|no uncertainty reported| 4427.60   A         | Broad-band measurement|189.497804 62.292517 (J2000)| Flux in fixed aperture|3" diameter aperture                    |Averaged from previously published data
3|V (HST/ACS) AB      | 22.514    ||mag                 |5.08E+14|  3.58E-06||Jy|2007ApJ...660...81M|no uncertainty reported|    5907   A         | Broad-band measurement|12 37 59.473 +62 17 33.06 (J2000)| Flux integrated from map|                                        |From reprocessed raw data; Corrected for contaminatingsources
4|R (Keck II) AB      | 22.74     || mag                |4.62E+14|  2.91E-06||Jy|2004AJ....127.3121W|no uncertainty reported|   648.7   A         | Broad-band measurement|12 37 59.473 +62 17 33.06 (J2000)| Total flux|                                        |From new raw data
5|R (Subaru) AB       | 22.64     ||mag                 |4.59E+14|  3.19E-06||Jy|2006ApJ...653.1027W|no uncertainty reported| 6534.16   A         | Broad-band measurement|189.497804 62.292517 (J2000)| Flux in fixed aperture|3" diameter aperture                    |Averaged from previously published data
6|i F775W (HST/ACS) AB      | 21.735    ||mag                 |3.86E+14|  7.35E-06||Jy|2007ApJ...660...81M|no uncertainty reported|    7764   A         | Broad-band measurement|12 37 59.473 +62 17 33.06 (J2000)| Flux integrated from map|                                        |From reprocessed raw data; Corrected for contaminatingsources
7|I (Subaru) AB       | 22.05     ||mag                 |3.76E+14|  5.50E-06||Jy|2006ApJ...653.1027W|no uncertainty reported| 7975.89   A         | Broad-band measurement|189.497804 62.292517 (J2000)| Flux in fixed aperture|3" diameter aperture                    |Averaged from previously published data
8|z F850LP (HST/ACS) AB      | 21.193    ||mag                 |3.17E+14|  1.21E-05||Jy|2007ApJ...660...81M|no uncertainty reported|    9445   A         | Broad-band measurement|12 37 59.473 +62 17 33.06 (J2000)| Flux integrated from map|                                        |From reprocessed raw data; Corrected for contaminatingsources
9|HK' (QUIRC) AB      | 20.48     |+/-0.15 |mag                 |1.58E+14|  2.33E-05|+/-3.22E-06|Jy|2006ApJ...653.1027W|uncertainty|18947.38   A         | Broad-band measurement|189.497804 62.292517 (J2000)| Flux in fixed aperture|3" diameter aperture                    |Averaged from previously published data
10|3.6 microns (IRAC)  | 41.60     |+/-2.08 |microJy             |8.44E+13|  4.16E-05|+/-2.08E-06|Jy|2011AJ....141....1T|rms uncertainty|     3.550 microns   | Broad-band measurement|189.497803 62.292522 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
11|4.5 microns (IRAC)  | 32.00     |+/-1.60 |microJy             |6.67E+13|  3.20E-05|+/-1.60E-06|Jy|2011AJ....141....1T|rms uncertainty|     4.493 microns   | Broad-band measurement|189.497803 62.292522 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
12|5.8 microns (IRAC)  | 23.30     |+/-1.26 |microJy             |5.23E+13|  2.33E-05|+/-1.26E-06|Jy|2011AJ....141....1T|rms uncertainty|     5.731 microns   | Broad-band measurement|189.497803 62.292522 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
13|8.0 microns (IRAC)  | 23.20     |+/-1.28 |microJy             |3.81E+13|  2.32E-05|+/-1.28E-06|Jy|2011AJ....141....1T|rms uncertainty|     7.872 microns   | Broad-band measurement|189.497803 62.292522 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
14|16 microns (IRS)    | 236.9     |+/-15.7 |microJy             |1.90E+13|  2.37E-04|+/-1.57E-05|Jy|2011AJ....141....1T|rms uncertainty|      15.8 microns   | Broad-band measurement|189.497803 62.292522 (J2000)| From fitting to map|                                        |From new raw data
15|24 microns (MIPS)   | 215.0     |+/-4.9  |microJy             |1.27E+13|  2.15E-04|+/-4.90E-06|Jy|2011AJ....141....1T|rms uncertainty|     23.68 microns   | Broad-band measurement|189.497803 62.292522 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
16|24 microns (MIPS)   | 221.5     |+/-2.6  |microJy             |1.27E+13|  2.21E-04|+/-2.60E-06|Jy|2011A&A...528A..35M|uncertainty|     23.68 microns   | Broad-band measurement|12 37 59.47 +62 17 33.01 (J2000)| Flux integrated from map|                                        |From new raw data
1|MIPS 24 microns     | 217.    |+/-7.0 |microJy         |1.25E+13 |  217.E-06|+/-7.0E-06|Jy |1990IRASF.C...0000M|3sigma uncertainty| 25        microns   | Broad-band measurement|115813.1 +302058 (B1950)| Flux in fixed aperture|                                        |From new raw data
17|70 microns (MIPS)   ||<4.4       |milliJy             |4.20E+12||4.40E-03|Jy|2011A&A...528A..35M|no uncertainty reported|     71.42 microns   | Broad-band measurement|12 37 59.47 +62 17 33.01 (J2000)| Flux integrated from map|                                        |From new raw data
2|70 microns (PACS)   |         |<2.4   |mJy             |4.283e+12|          |2.4E-03   |Jy |2.40e+01           |3sigma |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
3|100 microns (PACS)  | 1.2     |+/-0.4 |mJy             |2.998e+12|  1.2E-03 |+/-0.4E-03|Jy |2.40e+01           |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
4|160 microns (PACS)  | 5.3     |+/-1.7 |mJy             |1.874e+12|  5.3E-03 |+/-1.7E-03|Jy |2.40e+01           |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
5|250 microns (SPIRE) | 10.0    |+/-2.5 |mJy             |1.199e+12|  10.0E-03|+/-2.5e-03|Jy |2.40e+01           |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
6|350 microns (SPIRE) |         |<9.0   |mJy             |8.565e+11|          |9.0e-03   |Jy |2.40e+01           |3sigma |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
7|500 microns (SPIRE) |         |<12.0  |mJy             |5.996e+11|          |12.0e-03  |Jy |2.40e+01           |3sigma |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
8|1160 microns (Penner)|        |<2.1   |mJy             |2.58442E+11|        |2.1E-03   |Jy |2004MNRAS.354..779G|3sigma uncertainty|      1200 microns   | Broad-band measurement|16 36 55.9 +40 59 12 (J2000)| Flux integrated from map|S/N = 3.66                              |From new raw data
