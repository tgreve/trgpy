
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-02-19T11:09:36PST



Photometric Data for AzGN 15

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|4.0-8 keV (Chandra) | 1.11E-15  | |ergs cm^-2^ s^-1^   |1.45E+18|  7.65E-11| |Jy|2003AJ....126..539A|no uncertainty reported|       6   keV       | Broad-band measurement|12 35 49.44 +62 15 36.9 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
2|4-8 keV (Chandra)   | 0.91E-15  |+/-4   %|erg cm^-2^ s^-1^    |1.45E+18|  6.28E-11|+/-2.51E-12|Jy|2001AJ....122.2810B|estimated error|       6   keV       | Broad-band measurement|12 35 49.40 +62 15 36.8 (J2000)| Flux in fixed aperture|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
3|2-10 keV (Chandra)  | 1.20E-15  | |erg/cm^2^/s         |1.45E+18|  8.28E-11| |Jy|2009A&A...507..747G|no uncertainty reported|      6.00 keV       | Broad-band measurement|12 35 49.44 +62 15 36.9 (J2000)| Flux integrated from map|Observed flux                           |From new raw data; NED frequency assigned to mid-point ofband in keV
4|2-8 keV (Chandra)   | 1.02E-15  |+/-4   %|erg cm^-2^ s^-1^    |1.21E+18|  8.43E-11|+/-3.37E-12|Jy|2001AJ....122.2810B|estimated error|       5   keV       | Broad-band measurement|12 35 49.40 +62 15 36.8 (J2000)| Flux in fixed aperture|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
5|2.0-8 keV (Chandra) | 1.20E-15  | |ergs cm^-2^ s^-1^   |1.21E+18|  9.93E-11| |Jy|2003AJ....126..539A|no uncertainty reported|       5   keV       | Broad-band measurement|12 35 49.44 +62 15 36.9 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
6|0.5-8 keV (Chandra) | 1.20E-15  |+/-4   %|erg cm^-2^ s^-1^    |1.03E+18|  1.17E-10|+/-4.66E-12|Jy|2001AJ....122.2810B|estimated error|    4.25   keV       | Broad-band measurement|12 35 49.40 +62 15 36.8 (J2000)| Flux in fixed aperture|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
7|0.5-8 keV (Chandra) | 1.34E-15  | |ergs cm^-2^ s^-1^   |1.03E+18|  1.30E-10| |Jy|2003AJ....126..539A|no uncertainty reported|    4.25   keV       | Broad-band measurement|12 35 49.44 +62 15 36.9 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
8|2.0-4 keV (Chandra) | 0.25E-15  | |ergs cm^-2^ s^-1^   |7.25E+17|  3.45E-11| |Jy|2003AJ....126..539A|no uncertainty reported|       3   keV       | Broad-band measurement|12 35 49.44 +62 15 36.9 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
9|1.0-2 keV (Chandra) | 0.08E-15  | |ergs cm^-2^ s^-1^   |3.63E+17|  2.21E-11| |Jy|2003AJ....126..539A|no uncertainty reported|     1.5   keV       | Broad-band measurement|12 35 49.44 +62 15 36.9 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
10|0.5-2 keV (Chandra) | 0.12E-15  | |ergs cm^-2^ s^-1^   |3.02E+17|  3.97E-11| |Jy|2003AJ....126..539A|no uncertainty reported|    1.25   keV       | Broad-band measurement|12 35 49.44 +62 15 36.9 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
11|0.5-2 keV (Chandra) | 0.16E-15  |+/-4   %|erg cm^-2^ s^-1^    |3.02E+17|  5.30E-11|+/-2.12E-12|Jy|2001AJ....122.2810B|estimated error|    1.25   keV       | Broad-band measurement|12 35 49.40 +62 15 36.8 (J2000)| Flux in fixed aperture|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
12|0.5-1 keV (Chandra) | |<0.06E-15  |ergs cm^-2^ s^-1^   |1.81E+17| |3.31E-11|Jy|2003AJ....126..539A|3 sigma|    0.75   keV       | Broad-band measurement|12 35 49.44 +62 15 36.9 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
13|U (KPNO/MOSAIC) AB  | 24.61     |+/-0.10 |mag                 |8.44E+14|  5.20E-07|+/-4.79E-08|Jy|2005ApJ...635..853B|uncertainty|    3552   A         | Broad-band measurement|123549.44 +621536.8 (J2000)| Flux in fixed aperture|3" aperture                             |Averaged new and previously published data
14|[O II] 3727 (SUBARU)| 2.9E-16   |+/-0.8E-16|ergs cm^-2^ s^-1^   |8.04E+14|  3.61E-08|+/-9.95E-09|Jy|2006ApJ...651..713T|uncertainty|    3727   A         | Line measurement; flux integrated over line; lines measured in emission| | Flux integrated from map|                                        |From new raw data
15|B (SUBARU) AB       | 23.93     |+/-0.07 |mag                 |6.81E+14|  9.73E-07|+/-6.27E-08|Jy|2005ApJ...635..853B|uncertainty|    4400   A         | Broad-band measurement|123549.44 +621536.8 (J2000)| Flux in fixed aperture|3" aperture                             |Averaged new and previously published data
16|H{beta} (SUBARU)    | 1.6E-16   |+/-1.0E-16|ergs cm^-2^ s^-1^   |6.17E+14|  2.59E-08|+/-1.62E-08|Jy|2006ApJ...651..713T|uncertainty|    4861   A         | Line measurement; flux integrated over line; lines measured in emission| | Flux integrated from map|                                        |From new raw data
17|[O III] 4959 SUBARU | 1.9E-16   |+/-0.8E-16|ergs cm^-2^ s^-1^   |6.05E+14|  3.14E-08|+/-1.32E-08|Jy|2006ApJ...651..713T|uncertainty|    4959   A         | Line measurement; flux integrated over line; lines measured in emission| | Flux integrated from map|                                        |From new raw data
18|[O III] 5007 SUBARU | 6.4E-16   |+/-1.3E-16|ergs cm^-2^ s^-1^   |5.99E+14|  1.07E-07|+/-2.17E-08|Jy|2006ApJ...651..713T|uncertainty|    5007   A         | Line measurement; flux integrated over line; lines measured in emission| | Flux integrated from map|                                        |From new raw data
19|V (SUBARU) AB       | 23.60     |+/-0.04 |mag                 |5.42E+14|  1.32E-06|+/-4.86E-08|Jy|2005ApJ...635..853B|uncertainty|    5530   A         | Broad-band measurement|123549.44 +621536.8 (J2000)| Flux in fixed aperture|3" aperture                             |Averaged new and previously published data
20|R (SUBARU) AB       | 23.27     |+/-0.03 |mag                 |4.68E+14|  1.79E-06|+/-4.94E-08|Jy|2005ApJ...635..853B|uncertainty|    6400   A         | Broad-band measurement|123549.44 +621536.8 (J2000)| Flux in fixed aperture|3" aperture                             |Averaged new and previously published data
21|H{alpha} (SUBARU)   | 15.0E-16  |+/-1.0E-16|ergs cm^-2^ s^-1^   |4.57E+14|  3.28E-07|+/-2.19E-08|Jy|2006ApJ...651..713T|uncertainty|    6563   A         | Line measurement; flux integrated over line; lines measured in emission| | Flux integrated from map|                                        |From new raw data
22|I (SUBARU) AB       | 23.01     |+/-0.04 |mag                 |3.79E+14|  2.27E-06|+/-8.36E-08|Jy|2005ApJ...635..853B|uncertainty|    7900   A         | Broad-band measurement|123549.44 +621536.8 (J2000)| Flux in fixed aperture|3" aperture                             |Averaged new and previously published data
23|I (Cousins)         | 22.55     |+/-0.02 |mag                 |3.79E+14|  2.44E-06|+/-4.53E-08|Jy|2004ApJ...616...71S|1 sigma|    7900   A         | Broad-band measurement| | Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
24|z' (SUBARU) AB      | 22.84     |+/-0.05 |mag                 |3.30E+14|  2.65E-06|+/-1.22E-07|Jy|2005ApJ...635..853B|uncertainty|    9097   A         | Broad-band measurement|123549.44 +621536.8 (J2000)| Flux in fixed aperture|3" aperture                             |Averaged new and previously published data
3|HST F110W (WFC)      | 22.80     |+/-0.02 |mag             |2.67195e+14|  2.75423e-06|+/-5.0734774e-08|Jy |2011ApJ...728L...4H|uncertainty|     3.550 microns   | Broad-band measurement|09 03 11.6 +00 39 06 (J2000)| Flux in fixed aperture|                                        |From new raw data
25|J (Hale/WIRC) AB    | 21.77     |+/-0.07 |mag                 |2.40E+14|  7.11E-06|+/-4.59E-07|Jy|2005ApJ...635..853B|uncertainty|   1.250   microns   | Broad-band measurement|123549.44 +621536.8 (J2000)| Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
26|J (2MASS)           | 20.82     |+/-0.06 |mag                 |2.40E+14|  7.48E-06|+/-4.25E-07|Jy|2004ApJ...616...71S|1 sigma|    1.25   microns   | Broad-band measurement| | Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
6|F160W (HST/NICMOS)  | 21.92    |+/-0.01| mag                |1.87E+14|  6.19441e-06|+/-5.7052611e-08|Jy|2007A&A...470..467C|internal error|       1.6 microns   | Broad-band measurement| | From fitting to map|                                        |From new raw data
27|K_s_ (Hale/WIRC) AB | 21.49     |+/-0.18 |mag                 |1.39E+14|  9.21E-06|+/-1.53E-06|Jy|2005ApJ...635..853B|uncertainty|   2.150   microns   | Broad-band measurement|123549.44 +621536.8 (J2000)| Flux in fixed aperture|4" aperture; from 2004AJ....127..180C   |Averaged from previously published data
28|3.6 microns (IRAC)  | 3.4903E+01|+/-8.6256E-02|microJy             |8.44E+13|  3.49E-05|+/-8.63E-08|Jy|2013SSTSLC4.2....0C|uncertainty|3.55       microns   | Broad-band measurement|| Flux in fixed aperture|3.8" aperture                           |From new raw data
29|3.6 microns (IRAC)  | 4.2278E+01|+/-1.2167E-01|microJy             |8.44E+13|  4.23E-05|+/-1.22E-07|Jy|2013SSTSLC4.2....0C|uncertainty|3.55       microns   | Broad-band measurement|| Flux in fixed aperture|5.8" aperture                           |From new raw data
30|4.5 microns (IRAC)  | 4.4620E+01|+/-9.5700E-02|microJy             |6.67E+13|  4.46E-05|+/-9.57E-08|Jy|2013SSTSLC4.2....0C|uncertainty|4.493      microns   | Broad-band measurement|| Flux in fixed aperture|3.8" aperture                           |From new raw data
31|4.5 microns (IRAC)  | 5.2806E+01|+/-1.5404E-01|microJy             |6.67E+13|  5.28E-05|+/-1.54E-07|Jy|2013SSTSLC4.2....0C|uncertainty|4.493      microns   | Broad-band measurement|| Flux in fixed aperture|5.8" aperture                           |From new raw data
28|4.5 microns IRAC AB | 19.67     |+/-0.30 |mag                 |6.67E+13|  4.92E-05|+/-1.36E-05|Jy|2005ApJ...635..853B|uncertainty|   4.493   microns   | Broad-band measurement|123549.44 +621536.8 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged new and previously published data
29|4.5 microns (IRAC)  | 46.5      |+/-12.4 |microJy             |6.67E+13|  4.65E-05|+/-1.24E-05|Jy|2009ApJ...699.1610H|uncertainty|     4.493 microns   | Broad-band measurement|12 35 49.28 +62 15 36.5 (J2000)| Flux in fixed aperture|                                        |From new raw data
34|5.8 microns (IRAC)  | 6.2186E+01|+/-8.2192E-01|microJy             |5.23E+13|  6.22E-05|+/-8.22E-07|Jy|2013SSTSLC4.2....0C|uncertainty|5.731      microns   | Broad-band measurement|| Flux in fixed aperture|5.8" aperture                           |From new raw data
35|5.8 microns (IRAC)  | 5.8501E+01|+/-5.7076E-01|microJy             |5.23E+13|  5.85E-05|+/-5.71E-07|Jy|2013SSTSLC4.2....0C|uncertainty|5.731      microns   | Broad-band measurement|| Flux in fixed aperture|3.8" aperture                           |From new raw data
30|5.8 microns IRAC AB | 19.45     |+/-0.30 |mag                 |5.23E+13|  6.03E-05|+/-1.67E-05|Jy|2005ApJ...635..853B|uncertainty|   5.731   microns   | Broad-band measurement|123549.44 +621536.8 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged new and previously published data
31|5.8 microns (IRAC)  | 61.3      |+/-6.8  |microJy             |5.23E+13|  6.13E-05|+/-6.80E-06|Jy|2009ApJ...699.1610H|uncertainty|     5.731 microns   | Broad-band measurement|12 35 49.28 +62 15 36.5 (J2000)| Flux in fixed aperture|                                        |From new raw data
32|PAH 7.7 (Spitzer)   | 4.80E-15  |+/-0.65E-15|erg/s/cm^2^         |3.89E+13|  1.23E-05|+/-1.67E-06|Jy|2009ApJ...699..667M|rms uncertainty|       7.7 microns   | Line measurement; flux integrated over line; lines measured in emission|12 35 49.44 +62 15 36.8 (J2000)| Flux integrated from map|                                        |From new raw data
33|8.0 microns (IRAC)  | 64.1      |+/-22.0 |microJy             |3.85E+13|  6.41E-05|+/-2.20E-05|Jy|2009ApJ...699.1610H|uncertainty|     7.782 microns   | Broad-band measurement|12 35 49.28 +62 15 36.5 (J2000)| Flux in fixed aperture|                                        |From new raw data
34|8.0 microns IRAC AB | 19.36     |+/-0.30 |mag                 |3.81E+13|  6.55E-05|+/-1.81E-05|Jy|2005ApJ...635..853B|uncertainty|   7.872   microns   | Broad-band measurement|123549.44 +621536.8 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged new and previously published data
41|8.0 microns (IRAC)  | 6.3181E+01|+/-6.3401E-01|microJy             |3.81E+13|  6.32E-05|+/-6.34E-07|Jy|2013SSTSLC4.2....0C|uncertainty|7.872      microns   | Broad-band measurement|| Flux in fixed aperture|3.8" aperture                           |From new raw data
42|8.0 microns (IRAC)  | 7.2560E+01|+/-8.4855E-01|microJy             |3.81E+13|  7.26E-05|+/-8.49E-07|Jy|2013SSTSLC4.2....0C|uncertainty|7.872      microns   | Broad-band measurement|| Flux in fixed aperture|5.8" aperture                           |From new raw data
35|PAH 8.6 (Spitzer)   | 0.67E-15  |+/-0.07E-15|erg/s/cm^2^         |3.49E+13|  1.92E-06|+/-2.01E-07|Jy|2009ApJ...699..667M|rms uncertainty|       8.6 microns   | Line measurement; flux integrated over line; lines measured in emission|12 35 49.44 +62 15 36.8 (J2000)| Flux integrated from map|                                        |From new raw data
36|24 microns (MIPS)   | 585.6     | |microJy             |1.27E+13|  5.86E-04| |Jy|2007ApJ...660..167D|no uncertainty reported|   23.68   microns   | Broad-band measurement|12 35 49.43 +62 15 36.52 (J2000)| Flux in fixed aperture|                                        |From new raw data
37|24 microns (MIPS)   | 172.0     |+/-35.0 |microJy             |1.27E+13|  1.72E-04|+/-3.50E-05|Jy|2009ApJ...699.1610H|uncertainty|     23.68 microns   | Broad-band measurement|123549.44 +621536.8 (J2000)| Flux in fixed aperture|                                        |From new raw data
38|24 microns (Spitzer)| 630       | |microJy             |1.27E+13|  6.30E-04| |Jy|2011ApJ...726...93R|no uncertainty reported|     23.68 microns   | Broad-band measurement|12 35 49.44 +62 15 36.8 (J2000)| Not reported in paper|                                        |Averaged from previously published data
47|24 microns (MIPS)   | 6.4500E+02|+/-7.7617E+00|microJy             |1.27E+13|  6.45E-04|+/-7.76E-06|Jy|2013SSTSLC4.2....0C|uncertainty|23.68      microns   | Broad-band measurement|| Modelled datum|PSF fit                                 |From new raw data
48|24 microns (MIPS)   | 6.9596E+02|+/-6.8381E+00|microJy             |1.27E+13|  6.96E-04|+/-6.84E-06|Jy|2013SSTSLC4.2....0C|uncertainty|23.68      microns   | Broad-band measurement|| Flux in fixed aperture|14.7" aperture                          |From new raw data
39|70 microns (MIPS)   | |<4.1       |mJy             |4.20E+12| |4.10E-03|Jy|2009ApJ...699.1610H|3 sigma|     71.42 microns   | Broad-band measurement|123549.44 +621536.8 (J2000)| Flux in fixed aperture|                                        |From new raw data
40|CO 6-5 line (PdBI)  | 2.3       |+/-0.4  |Jy km s^-1^         |6.91E+11|  7.49E-07|+/-1.30E-07|Jy|2006ApJ...640..228T|uncertainty|   2.202             | Line measurement; flux integrated over line; lines measured in emission|12 35 49.42 +62 15 36.9 (J2000)| Flux integrated from map|                                        |From new raw data
41|850 microns (SCUBA) | 8.3       |+/-2.5  |milliJy             |3.53E+11|  8.30E-03|+/-2.50E-03|Jy|2005ApJ...622..772C|uncertainty|     850   microns   | Broad-band measurement|123549.44 +621536.8 (J2000)| Flux integrated from map|                                        |From new raw data
42|CO 3-2 line (PdBI)  | 1.6       |+/-0.2  |Jy km s^-1^         |3.46E+11|  5.20E-07|+/-6.50E-08|Jy|2006ApJ...640..228T|uncertainty|   2.202             | Line measurement; flux integrated over line; lines measured in emission|12 35 49.42 +62 15 36.9 (J2000)| Flux integrated from map|                                        |From new raw data
43|1.3 mm (PdBI)       | 2.0       |+/-0.6  |milliJy             |2.31E+11|  2.00E-03|+/-6.00E-04|Jy|2006ApJ...640..228T|uncertainty|     1.3   mm        | Broad-band measurement| | Flux integrated from map|                                        |From new raw data
44|1.4 GHz (VLA)       | 104       |+/-8    | microJy            |1.40E+09|  1.04E-04|+/-8.00E-06|Jy|2006MNRAS.371..963B|1 sigma|       1.4 GHz       | Broad-band measurement|12 35 49.431 +62 15 36.71 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
45|1.4 GHz (VLA)       | 93.1      |+/-6.4  |microJy             |1.40E+09|  9.31E-05|+/-6.40E-06|Jy|2010ApJS..188..178M|uncertainty|       1.4 GHz       | Broad-band measurement|12 35 49.41 +62 15 36.9 (J2000)| Total flux; Beam filling or dilution corrected|Major=0.9"; Minor=0.0"; PA=140 deg      |From new raw data
46|1.4 GHz (VLA)       | 74.6      |+/-9.5  |microJy             |1.40E+09|  7.46E-05|+/-9.50E-06|Jy|2000ApJ...533..611R|1 sigma|1.4        GHz       | Broad-band measurement; broad-band flux derived by integration over spectrum; synthetic band|123549.438 +621536.75 (J2000)| Flux integrated from map; Pointing and beam filling|                                        |From new raw data; Corrected for contaminating sources
