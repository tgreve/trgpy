
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-03-28T04:53:10PDT



Photometric Data for CFRS 03.0346

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|F450W (HST)         | 23.77     | | mag                |6.63E+14|  1.35E-06| |Jy|2004A&A...421..847Z|no uncertainty reported|    4519   A         | Broad-band measurement| | Flux in fixed aperture|3" aperture                             |From reprocessed raw data
2|H{beta} (VLT)       | 1.9E-16   |+/-1.1E-16|ergs cm^-2^ s^-1^   |6.17E+14|  3.08E-08|+/-1.78E-08|Jy|2006ApJ...651..713T|uncertainty|    4861   A         | Line measurement; flux integrated over line; lines measured in emission| | Flux integrated from map|                                        |From new raw data
3|[O III] 4959 (VLT)  | 7.2E-16   |+/-2.6E-16|ergs cm^-2^ s^-1^   |6.05E+14|  1.19E-07|+/-4.30E-08|Jy|2006ApJ...651..713T|uncertainty|    4959   A         | Line measurement; flux integrated over line; lines measured in emission| | Flux integrated from map|                                        |From new raw data
4|[O III] 5007 (VLT)  | 10.7E-16  |+/-3.2E-16|ergs cm^-2^ s^-1^   |5.99E+14|  1.79E-07|+/-5.34E-08|Jy|2006ApJ...651..713T|uncertainty|    5007   A         | Line measurement; flux integrated over line; lines measured in emission| | Flux integrated from map|                                        |From new raw data
5|H{alpha} (VLT)      | 15.2E-16  |+/-2.0E-16|ergs cm^-2^ s^-1^   |4.57E+14|  3.33E-07|+/-4.38E-08|Jy|2006ApJ...651..713T|uncertainty|    6563   A         | Line measurement; flux integrated over line; lines measured in emission| | Flux integrated from map|                                        |From new raw data
6|I (Cousins)         | 21.29     |+/-0.05 |mag                 |3.79E+14|  7.77E-06|+/-3.66E-07|Jy|2004ApJ...616...71S|1 sigma|    7900   A         | Broad-band measurement| | Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
7|F814W (HST)         | 21.52     | | mag                |3.78E+14|  6.14E-06| |Jy|2004A&A...421..847Z|no uncertainty reported|    7924   A         | Broad-band measurement| | Flux in fixed aperture|3" aperture                             |From reprocessed raw data
8|J (2MASS)           | 19.66     |+/-0.04 |mag                 |2.40E+14|  2.18E-05|+/-8.17E-07|Jy|2004ApJ...616...71S|1 sigma|    1.25   microns   | Broad-band measurement| | Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
9|F160W (HST) AB      | 20.73     |+/-0.02 |mag                 |1.87E+14|  1.85E-05|+/-3.41E-07|Jy|2010MNRAS.405..234S|uncertainty|      1.60 microns   | Broad-band measurement|03 02 27.73 +00 06 53.5 (J2000)| Flux in fixed aperture|                                        |From new raw data
10|K_s_ (2MASS)        | 19.14     |+/-0.03 |mag                 |1.38E+14|  1.47E-05|+/-4.13E-07|Jy|2004ApJ...616...71S|1 sigma|    2.17   microns   | Broad-band measurement| | Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
11|K (UKIRT)           | 18.33     |+/-0.02 | mag                |1.36E+14|  3.06E-05|+/-5.63E-07|Jy|2004MNRAS.351..447C|uncertainty|     2.2   microns   | Broad-band measurement|03 02 27.72 +00 06 53.2 (J2000)| Flux in fixed aperture|3" diameter aperture                    |From new raw data
12|3.6 microns (IRAC)  | 75.8      |+/-7.7  |microJy             |8.44E+13|  7.58E-05|+/-7.70E-06|Jy|2009ApJ...699.1610H|uncertainty|     3.550 microns   | Broad-band measurement|03 02 27.74 +00 06 53.4 (J2000)| Flux in fixed aperture|                                        |From new raw data
13|4.5 microns (IRAC)  | 81.6      |+/-8.3  |microJy             |6.67E+13|  8.16E-05|+/-8.30E-06|Jy|2009ApJ...699.1610H|uncertainty|     4.493 microns   | Broad-band measurement|03 02 27.74 +00 06 53.4 (J2000)| Flux in fixed aperture|                                        |From new raw data
14|5.8 microns (IRAC)  | 61.5      |+/-6.5  |microJy             |5.23E+13|  6.15E-05|+/-6.50E-06|Jy|2009ApJ...699.1610H|uncertainty|     5.731 microns   | Broad-band measurement|03 02 27.74 +00 06 53.4 (J2000)| Flux in fixed aperture|                                        |From new raw data
15|PAH 6.2 (Spitzer)   | 2.29E-15  |+/-0.46E-15|erg/s/cm^2^         |4.84E+13|  4.73E-06|+/-9.50E-07|Jy|2009ApJ...699..667M|rms uncertainty|       6.2 microns   | Line measurement; flux integrated over line; lines measured in emission|03 02 27.73 +00 06 53.5 (J2000)| Flux integrated from map|                                        |From new raw data
16|PAH 7.7 (Spitzer)   | 8.49E-15  |+/-1.05E-15|erg/s/cm^2^         |3.89E+13|  2.18E-05|+/-2.70E-06|Jy|2009ApJ...699..667M|rms uncertainty|       7.7 microns   | Line measurement; flux integrated over line; lines measured in emission|03 02 27.73 +00 06 53.5 (J2000)| Flux integrated from map|                                        |From new raw data
17|8.0 microns (IRAC)  | 63.4      |+/-6.8  |microJy             |3.85E+13|  6.34E-05|+/-6.80E-06|Jy|2009ApJ...699.1610H|uncertainty|     7.782 microns   | Broad-band measurement|03 02 27.74 +00 06 53.4 (J2000)| Flux in fixed aperture|                                        |From new raw data
18|PAH 8.6 (Spitzer)   | 3.29E-15  |+/-0.67E-15|erg/s/cm^2^         |3.49E+13|  9.43E-06|+/-1.92E-06|Jy|2009ApJ...699..667M|rms uncertainty|       8.6 microns   | Line measurement; flux integrated over line; lines measured in emission|03 02 27.73 +00 06 53.5 (J2000)| Flux integrated from map|                                        |From new raw data
19|PAH 11.3 (Spitzer)  | 2.27E-15  |+/-0.47E-15|erg/s/cm^2^         |2.65E+13|  8.57E-06|+/-1.77E-06|Jy|2009ApJ...699..667M|rms uncertainty|      11.3 microns   | Line measurement; flux integrated over line; lines measured in emission|03 02 27.73 +00 06 53.5 (J2000)| Flux integrated from map|                                        |From new raw data
20|PAH 12.7 (Spitzer)  | 2.88E-15  |+/-0.45E-15|erg/s/cm^2^         |2.36E+13|  1.22E-05|+/-1.91E-06|Jy|2009ApJ...699..667M|rms uncertainty|      12.7 microns   | Line measurement; flux integrated over line; lines measured in emission|03 02 27.73 +00 06 53.5 (J2000)| Flux integrated from map|                                        |From new raw data
21|15 microns (ISO)    | 254       |+/-96   |microJy             |2.00E+13|  2.54E-04|+/-9.60E-05|Jy|2003ApJ...587...41W|uncertainty|    15.0   microns   | Broad-band measurement| | Flux in fixed aperture|                                        |From new raw data
22|24 microns (MIPS)   | 0.23      |+/-10  %|milliJy             |1.27E+13|  2.30E-04|+/-2.30E-05|Jy|2009A&A...502..541E|uncertainty|     23.68 microns   | Broad-band measurement| | Flux in fixed aperture|                                        |From reprocessed raw data
23|24 microns (MIPS)   | 479.0     |+/-53.0 |microJy             |1.27E+13|  4.79E-04|+/-5.30E-05|Jy|2009ApJ...699.1610H|uncertainty|     23.68 microns   | Broad-band measurement|030227.73 +000653.5 (J2000)| Flux in fixed aperture|                                        |From new raw data
24|70 microns (MIPS)   | |<8.8       |milliJy             |4.20E+12| |8.80E-03|Jy|2009A&A...502..541E|3 sigma|     71.42 microns   | Broad-band measurement| | Flux in fixed aperture|                                        |From reprocessed raw data
25|70 microns (MIPS)   | |<13.6      |milliJy             |4.20E+12| |1.36E-02|Jy|2009ApJ...699.1610H|3 sigma|     71.42 microns   | Broad-band measurement|030227.73 +000653.5 (J2000)| Flux in fixed aperture|                                        |From new raw data
26|350 microns (SHARC2)| 42.2      |+/-9.8  |milliJy             |8.57E+11|  4.22E-02|+/-9.80E-03|Jy|2006ApJ...650..592K|uncertainty|     350   microns   | Broad-band measurement| | Total flux|                                        |From new raw data
27|450 microns (SCUBA) | |<63        |milliJy             |6.66E+11| |6.30E-02|Jy|2003ApJ...587...41W|3 sigma|     450   microns   | Broad-band measurement|03 02 27.60 +00 06 52.5 (J2000)| Flux in fixed aperture|12" diameter aperture; S/N = 3.5        |From new raw data
28|850 microns (SCUBA) | 4.4       |+/-1.3  |milliJy             |3.53E+11|  4.40E-03|+/-1.30E-03|Jy|2005ApJ...622..772C|uncertainty|     850   microns   | Broad-band measurement|030227.73 +000653.5 (J2000)| Flux integrated from map|                                        |From new raw data
29|850 microns (SCUBA) | 4.4       |+/-1.3  |milliJy             |3.53E+11|  4.40E-03|+/-1.30E-03|Jy|2003ApJ...587...41W|uncertainty|     850   microns   | Broad-band measurement|03 02 27.60 +00 06 52.5 (J2000)| Flux in fixed aperture|12" diameter aperture; S/N = 3.5        |From new raw data
30|1.4 GHz (VLA)       | 226       |+/-12   |microJy             |1.40E+09|  2.26E-04|+/-1.20E-05|Jy|2003ApJ...587...41W|uncertainty|     1.4   GHz       | Broad-band measurement| | Peak flux|                                        |From new raw data
31|1.4 GHz (VLA)       | 226       |+/-12   | microJy            |1.40E+09|  2.26E-04|+/-1.20E-05|Jy|2004MNRAS.351..447C|uncertainty|     1.4   GHz       | Broad-band measurement|03 02 27.73 +00 06 53.5 (J2000)| Flux integrated from map|                                        |From new raw data
