

Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.


queryDateTime:2009-11-03T15:07:35PST



Photometric Data for HS1700.850.1 (z=2.816)




No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|U (WHT)             |       |>27.1  |mag                 |8.48549e+14|  |5.24809e-08|Jy|2004ApJ...616...71S|3sigma uncertainty|    1.25   microns   | Broad-band measurement| | Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
1|g (WHT)             | 27.0      |+/-0.3  |mag                 |6.17874e+14|5.75440e-08|+/-1.83136e-08 |Jy|2004ApJ...616...71S|sigma uncertainty|    1.25   microns   | Broad-band measurement| | Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
2|WHT/PPC Ra          | 26.1      |+/-0.3  |ABmag               |4.70E+14|  1.36E-07 |+/-0.43E-07|Jy|2004A&A...421..847Z|no uncertainty reported|    7924   A         | Broad-band measurement| | Flux in fixed aperture|3" aperture                             |From reprocessed raw data
3|HST/ACS F814W       | 25.8      |+/-0.2  |ABmag               |3.78E+14|  1.79E-07 |+/-0.36E-07|Jy|2004A&A...421..847Z|no uncertainty reported|    7924   A         | Broad-band measurement| | Flux in fixed aperture|3" aperture                             |From reprocessed raw data
4|P200/WIRC J         | 24.4      |+/-0.2  |ABmag               |2.40e+14|  6.49E-07 |+/-1.31E-07|Jy|2004A&A...421..847Z|no uncertainty reported|    7924   A         | Broad-band measurement| | Flux in fixed aperture|3" aperture                             |From reprocessed raw data
5|P200/WIRC Ks        | 23.20     |+/-0.13 |ABmag               |1.38e+14|  1.96E-06 |+/-0.25E-06|Jy|2004A&A...421..847Z|no uncertainty reported|    7924   A         | Broad-band measurement| | Flux in fixed aperture|3" aperture                             |From reprocessed raw data
6|IRAC 4.5um          | 10.2      |+/-0.9  |microJy             |6.67E+13|  10.2E-06 |+/-0.9E-06 |Jy|1996AJ....111.1431B|uncertainty|1.49       GHz       | Broad-band measurement| | Peak flux|                                        |From new raw data
7|IRAC 4.5um          | 10.2      |+/-0.9  |microJy             |6.67E+13|  10.2E-06 |+/-0.9E-06 |Jy|1996AJ....111.1431B|uncertainty|1.49       GHz       | Broad-band measurement| | Peak flux|                                        |From new raw data
8|IRAC 8um            | 13.2      |+/-1.2  |microJy             |3.81E+13|  13.2E-06 |+/-1.2E-06 |Jy|1996AJ....111.1431B|uncertainty|1.49       GHz       | Broad-band measurement| | Peak flux|                                        |From new raw data
9|MIPS 24um           | 171.0     |+/-7.0  |microJy             |1.27E+13|  171.0E-06|+/-7.0E-06 |Jy|1996AJ....111.1431B|uncertainty|1.49       GHz       | Broad-band measurement| | Peak flux|                                        |From new raw data
10|SCUBA-2 450um      | 45.0      |+/-6.0  |milliJy             |666.0E+09|  45.0E-03|+/-6.0E-03 |Jy|1996AJ....111.1431B|uncertainty|1.49       GHz       | Broad-band measurement| | Peak flux|                                        |From new raw data
11|SCUBA-2 850um      | 19.1      |+/-0.8  |milliJy             |353.0E+09|  19.1E-03|+/-0.8E-03 |Jy|1996AJ....111.1431B|uncertainty|1.49       GHz       | Broad-band measurement| | Peak flux|                                        |From new raw data
12|SMA 870um          | 14.5      |+/-1.1  |milliJy             |3.44589e+11|14.5E-03|+/-0.8E-03 |Jy|1996AJ....111.1431B|uncertainty|1.49       GHz       | Broad-band measurement| | Peak flux|                                        |From new raw data
13|IRAM PdBI 149.2GHz | 1.39      |+/-0.15 |milliJy             |149.2E+09|  1.39E-03|+/-0.15E-03|Jy|1996AJ....111.1431B|uncertainty|1.49       GHz       | Broad-band measurement| | Peak flux|                                        |From new raw data
14|IRAM PdBI 103.8GHz | 0.38      |+/-0.08 |milliJy             |103.8E+09|  0.38E-03|+/-0.08E-03|Jy|1996AJ....111.1431B|uncertainty|1.49       GHz       | Broad-band measurement| | Peak flux|                                        |From new raw data
15|IRAM PdBI 100.8GHz | 0.31      |+/-0.13 |milliJy             |100.8E+09|  0.31E-03|+/-0.13E-03|Jy|1996AJ....111.1431B|uncertainty|1.49       GHz       | Broad-band measurement| | Peak flux|                                        |From new raw data
16|IRAM PdBI 91.7GHz  | 0.25      |+/-0.07 |milliJy             |91.7E+09 |  0.25E-03|+/-0.07E-03|Jy|1996AJ....111.1431B|uncertainty|1.49       GHz       | Broad-band measurement| | Peak flux|                                        |From new raw data
