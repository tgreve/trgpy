
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-06-16T05:11:03PDT



Photometric Data for SDSS J142005.35+530115.4

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
5|K_s (PALOMAR DEEP2) VEGA     | 17.27     || mag                |1.39E+14|  7.66E-05||Jy|2007MNRAS.382..109T|no uncertainty reported|      2.15 microns   | Broad-band measurement|215.02251 +53.02097 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
6|24 microns (MIPS)   | 571.3     ||microJy             |1.27E+13|  5.71E-04||Jy|2011ApJ...726...93R|no uncertainty reported|     23.68 microns   | Broad-band measurement|14 20 05.43 +53 01 15.5 (J2000)| Not reported in paper|                                        |Averaged from previously published data
