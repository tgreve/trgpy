
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-07-08T06:53:30PDT



Photometric Data for SDSS J123707.83+621057.6

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|U (KPNO) AB         | 24.22     ||mag                 |8.44E+14|  7.45E-07||Jy|2006ApJ...653.1004R|no uncertainty reported|    3550   A         | Broad-band measurement|123707.82 +621057.6 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data; derived from aflux in a different band and a color
2|u (SDSS PSF) AB     | 23.671    |+/-0.737|asinh mag           |8.36E+14|  1.06E-06|+/-1.02E-06|Jy|2007SDSS6.C...0000:|based on count statistics only|3585       A         | Broad-band measurement|189.2826524315 62.1826913248 (J2000)| Modelled datum|SDSS flags: CANONICAL_CENTER - used canonical, not local, center; CHILD - object is part of a blended parent object; INTERP - object contains interpolated-over pixels; ELLIPFAINT - no isophotal fits performed; AMOMENT_FAINT - too faint for adaptive moments;|From new raw data
3|G (KECK) AB         | 23.67     ||mag                 |6.27E+14|  1.24E-06||Jy|2006ApJ...653.1004R|no uncertainty reported|    4780   A         | Broad-band measurement|123707.82 +621057.6 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data; derived from aflux in a different band and a color
4|g (SDSS PSF) AB     | 23.746    |+/-0.354|asinh mag           |6.17E+14|  1.06E-06|+/-4.06E-07|Jy|2007SDSS6.C...0000:|based on count statistics only|4858       A         | Broad-band measurement|189.2826524315 62.1826913248 (J2000)| Modelled datum|SDSS flags: CANONICAL_CENTER - used canonical, not local, center; CHILD - object is part of a blended parent object; NOPETRO - no Petrosian radius could be determined; PETROFAINT - Petrosian radius measured at very low surface brightness; ELLIPFAINT - no isophotal fits performed; AMOMENT_FAINT - too faint for adaptive moments;|From new raw data
5|r (SDSS PSF) AB     | 22.468    |+/-0.175|asinh mag           |4.77E+14|  3.69E-06|+/-6.11E-07|Jy|2007SDSS6.C...0000:|based on count statistics only|6290       A         | Broad-band measurement|189.2826524315 62.1826913248 (J2000)| Modelled datum|SDSS flags: CHILD - object is part of a blended parent object; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding; CANONICAL_BAND - this band was primary (usually r);|From new raw data
6|R (Keck II) AB      | 23.38     || mag                |4.62E+14|  1.61E-06||Jy|2004AJ....127.3121W|no uncertainty reported|   648.7   A         | Broad-band measurement|12 37 07.837 +62 10 57.65 (J2000)| Total flux|                                        |From new raw data
7|R (KECK) AB         | 23.16     ||mag                 |4.39E+14|  1.98E-06||Jy|2006ApJ...653.1004R|no uncertainty reported|    6830   A         | Broad-band measurement|123707.82 +621057.6 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data
8|i (SDSS PSF) AB     | 23.388    |+/-0.341|asinh mag           |3.89E+14|  1.34E-06|+/-5.87E-07|Jy|2007SDSS6.C...0000:|based on count statistics only|7706       A         | Broad-band measurement|189.2826524315 62.1826913248 (J2000)| Modelled datum|SDSS flags: CANONICAL_CENTER - used canonical, not local, center; CHILD - object is part of a blended parent object; MANYPETRO - more than one Petrosian radius; COSMIC_RAY - contains a cosmic ray pixel; INTERP - object contains interpolated-over pixels; PETROFAINT - Petrosian radius measured at very low surface brightness; ELLIPFAINT - no isophotal fits performed; AMOMENT_FAINT - too faint for adaptive moments;|From new raw data
9|z (SDSS PSF) AB     | 22.521    |+/-0.875|asinh mag           |3.25E+14|  1.51E-06|+/-4.42E-06|Jy|2007SDSS6.C...0000:|based on count statistics only|9222       A         | Broad-band measurement|189.2826524315 62.1826913248 (J2000)| Modelled datum|SDSS flags: CANONICAL_CENTER - used canonical, not local, center; CHILD - object is part of a blended parent object; MANYR50 - more than one 50% radius; MANYR90 - more than one 90% radius; ELLIPFAINT - no isophotal fits performed; AMOMENT_FAINT - too faint for adaptive moments;|From new raw data
10|J (WIRC) AB         | 22.02     ||mag                 |2.40E+14|  5.65E-06||Jy|2006ApJ...653.1004R|no uncertainty reported|   1.250   microns   | Broad-band measurement|123707.82 +621057.6 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data
11|K_s (WIRC) AB       | 21.47     ||mag                 |1.39E+14|  9.38E-06||Jy|2006ApJ...653.1004R|no uncertainty reported|   2.150   microns   | Broad-band measurement|123707.82 +621057.6 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data
12|3.6 microns IRAC AB | 21.15     |+/-0.07 |mag                 |8.44E+13|  1.26E-05|+/-8.12E-07|Jy|2006ApJ...653.1004R|uncertainty|   3.550   microns   | Broad-band measurement|123707.82 +621057.6 (J2000)| Flux integrated from map|                                        |From new raw data
13|4.5 microns IRAC AB | 21.05     |+/-0.07 |mag                 |6.67E+13|  1.38E-05|+/-8.90E-07|Jy|2006ApJ...653.1004R|uncertainty|   4.493   microns   | Broad-band measurement|123707.82 +621057.6 (J2000)| Flux integrated from map|                                        |From new raw data
14|5.8 microns IRAC AB | 21.19     |+/-0.17 |mag                 |5.23E+13|  1.21E-05|+/-1.90E-06|Jy|2006ApJ...653.1004R|uncertainty|   5.731   microns   | Broad-band measurement|123707.82 +621057.6 (J2000)| Flux integrated from map|                                        |From new raw data
15|24 microns (MIPS)   | 70.3      |+/-9.8  |microJy             |1.27E+13|  7.03E-05|+/-9.80E-06|Jy|2011A&A...528A..35M|uncertainty|     23.68 microns   | Broad-band measurement|12 37 07.83 +62 10 57.72 (J2000)| Flux integrated from map|                                        |From new raw data
1|24 microns (MIPS)   | 588       |+/-63   |mJy             |1.27E+13|588.E-03|+/-63.0E-03|Jy|2009ApJ...694.1517D|3sigma uncertainty|     23.68 microns   | Broad-band measurement|12 37 11.89 +62 22 11.8 (J2000)| Flux integrated from map|                                        |From new raw data
16|70 microns (MIPS)   ||<3.4       |milliJy             |4.20E+12||3.40E-03|Jy|2011A&A...528A..35M|no uncertainty reported|     71.42 microns   | Broad-band measurement|12 37 07.83 +62 10 57.72 (J2000)| Flux integrated from map|                                        |From new raw data
2|70 microns (MIPS)   |           |<2.6  |mJy             |4.20E+12| |2.6E-03|Jy|2009ApJ...699.1610H|3 sigma|     71.42 microns   | Broad-band measurement|221804.42 +002154.4 (J2000)| Flux in fixed aperture|                                        |From new raw data
3|850 microns (SCUBA) |           |<4.8    |mJy             |3.53E+11|  |4.8E-03|Jy|2005MNRAS.358..149P|3sigma uncertainty|     850   microns   | Broad-band measurement|12 37 11.7 +62 22 12 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
4|1200 microns (MAMBO)|           |<2.6    |mJy             |2.50E+11|        |2.6E-03|Jy|2004MNRAS.354..779G|3sigma uncertainty|      1200 microns   | Broad-band measurement|16 36 55.9 +40 59 12 (J2000)| Flux integrated from map|S/N = 3.66                              |From new raw data
5|1.4 GHz (VLA)       | 24.1     |+/-8.6  | microJy        |1.40E+09| 24.1E-06|+/-8.6E-06|Jy|2006MNRAS.371..963B|1 sigma|       1.4 GHz       | Broad-band measurement|16 36 55.767 +40 59 09.97 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
