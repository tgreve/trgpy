
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-07-10T13:42:15PDT



Photometric Data for SPT0551-50

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
5|250 microns (SPIRE)|  632.6   |+/-11.9 |mJy                 |1.199e+12| 632.6E-03|+/-11.9e-03 |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
6|350 microns (SPIRE)|  600.2   |+/-19.9  |mJy                |8.565e+11|600.2E-03 |+/-19.9e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
8|500 microns (SPIRE) | 420.3   |+/-11.9 |mJy                 |5.996e+11|420.3E-03 |+/-11.9e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
1|870 microns (LABOCA)| 138.7   |+/-4.4  |milliJy            |3.45E+11|  138.7E-03|+/-4.4E-03|Jy|2009ApJ...707.1201W|uncertainty|       870 microns   | Broad-band measurement|03 32 29.33 -27 56 19.3 (J2000)| Flux integrated from map|S/N = 4.6                               |From new raw data
1|1.4 mm (SPT)        | 35.9    |+/-6.8 |milliJy             |2.20E+11|  35.9E-03|+/-6.8E-03|Jy|2010ApJ...719..763V|uncertainty|       1.4 mm        | Broad-band measurement|74.804 -59.708 (J2000)| Flux integrated from map|De-boosted flux; S/N = 7.05             |From new raw data
3|2.0 mm (SPT)        | 10.5    |+/-1.6 |milliJy             |1.50E+11|  10.5E-03|+/-1.6E-03|Jy|2010ApJ...719..763V|uncertainty|       2.0 mm        | Broad-band measurement|74.804 -59.708 (J2000)| Flux integrated from map|De-boosted flux; S/N = 6.20             |From new raw data
