
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-05-28T01:42:09PDT



Photometric Data for HXMM01

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|NUV GALEX           |          |<0.5     |uJy |1.30E+15 |           |0.5E-06      |Jy|2011ApJ...728L...4H|3sigma uncertainty       | | | | |
2|u CFHT              | 0.5      |+/-0.1   |uJy |7.889E+14|0.5E-06    |+/-0.1E-06   |Jy|2011ApJ...728L...4H|uncertainty       | | | | |
3|g CFHT              | 1.3      |+/-0.1   |uJy |6.118E+14|1.3E-06    |+/-0.1E-06   |Jy|2011ApJ...728L...4H|uncertainty       | | | | |
4|r CFHT              | 2.3      |+/-0.2   |uJy |4.835E+14|2.3E-06    |+/-0.2E-06   |Jy|2011ApJ...728L...4H|uncertainty       | | | | |
5|i CFHT              | 2.5      |+/-0.3   |uJy |3.945E+14|2.5E-06    |+/-0.3E-06   |Jy|2011ApJ...728L...4H|uncertainty       | | | | |
6|z CFHT              | 3.8      |+/-0.6   |uJy |3.407E+14|3.8E-06    |+/-0.6E-06   |Jy|2011ApJ...728L...4H|uncertainty       | | | | |
7|F110W HST           | 6.2      |+/-0.4   |uJy |2.67195E+14|6.2E-06  |+/-0.4E-06   |Jy|2011ApJ...728L...4H|uncertainty       | | | | |
8|J WHT               | 6.8      |+/-0.8   |uJy |2.398E+14|6.8E-06    |+/-0.8E-06   |Jy|2011ApJ...728L...4H|uncertainty       | | | | |
9|K WHT               | 22.5     |+/-3.4   |uJy |1.394E+14|22.5E-06   |+/-3.4E-06   |Jy|2011ApJ...728L...4H|uncertainty       | | | | |
10|3.6 microns (IRAC) | 48.5     |+/-5.8   |uJy |8.44E+13 |48.5E-06   |+/-5.8E-06   |Jy|2011ApJ...728L...4H|uncertainty       | | | | |
11|4.5 microns (IRAC) | 64.1     |+/-5.9   |uJy |6.67E+13 |64.1E-06   |+/-5.9E-06   |Jy|2011ApJ...728L...4H|uncertainty       | | | | |
12|5.8 microns (IRAC) | 111.9    |+/-12.0  |uJy |5.23E+13 |111.9E-06  |+/-12.0E-06  |Jy|2009AJ....137.3884R|uncertainty       | | | | |
13|8.0 microns (IRAC) | 86.9     |+/-12.7  |uJy |3.85E+13 |86.9E-06   |+/-12.7E-06  |Jy|2009ApJ...699.1610H|uncertainty       | | | | |
14|24 microns (MIPS)  | 2280.    |+/-100.0 |uJy |1.27E+13 |2280.E-06  |+/-100.0E-06 |Jy|1990IRASF.C...0000M|3sigma uncertainty| | | | |
15|70 microns (PACS)  | 7970.    |+/-3890  |uJy |4.28e+12 |7970.E-06  |+/-3890.E-06 |Jy|Reference          |uncertainty       | | | | |
16|100 microns (PACS) | 31700.   |+/-3000  |uJy |2.998e+12|31700E-06  |+/-3000.E-06 |Jy|Reference          |uncertainty       | | | | |
17|160 microns (PACS) | 102100.  |+/-6000  |uJy |1.874e+12|102100.E-06|+/-6000.E-06 |Jy|Reference          |uncertainty       | | | | |
18|250 microns (SPIRE)| 180.3    |+/-14.3  |mJy |1.199e+12|180.3E-03  |+/-14.3E-03  |Jy|Reference          |uncertainty       | | | | |
19|350 microns (SPIRE)| 192.1    |+/-15.5  |mJy |8.57e+11|192.1E-03  |+/-15.5E-03  |Jy|Reference          |uncertainty       | | | | |
20|500 microns (SPIRE)| 131.6    |+/-11.3  |mJy |5.996e+11|131.6E-03  |+/-11.3E-03  |Jy|Reference          |uncertainty       | | | | |
21|880 microns (SMA)  | 27.0     |+/-3.0   |mJy |3.40673e+11|27.0E-03   |+/-3.00E-03  |Jy|2010ApJ...709..210K|uncertainty       | | | | |
22|1.2 mm (MAMBO)     | 11.2     |+/-1.9   |mJy |2.50E+11 |11.2E-03   |+/-1.9E-03   |Jy|2010A&A...522L...4L|uncertainty       | | | | |
23|2.1 mm (PdBI)      | 1.22     |+/-0.24  |mJy |1.43E+11 |1.22E-03   |+/-0.24E-03  |Jy|2010Natur.464..733S|uncertainty       | | | | |
24|1.4 GHz (VLA)      |          |<420.    |uJy |1.40E+09 |           |420.E-06|Jy|2007MNRAS.380..199I|3rms uncertainty|       1.4 GHz       | Broad-band measurement|10 52 28.995 +57 22 22.42 (J2000)| Flux integrated from map|                                        |From reprocessed raw data
