
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-07-10T12:46:28PDT



Photometric Data for PKS 0324-228

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|3.6 microns (IRAC)  | 39.4      |+/-4.2  | microJy            |8.44E+13|  3.94E-05|+/-4.20E-06|Jy|2007ApJS..171..353S|uncertainty|   3.550   microns   | Broad-band measurement|03 27 04.4 -22 39 42.60 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
2|4.5 microns (IRAC)  | 39.7      |+/-4.3  | microJy            |6.67E+13|  3.97E-05|+/-4.30E-06|Jy|2007ApJS..171..353S|uncertainty|   4.493   microns   | Broad-band measurement|03 27 04.4 -22 39 42.60 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
3|5.8 microns (IRAC)  | 61.1      |+/-8.6  | microJy            |5.23E+13|  6.11E-05|+/-8.60E-06|Jy|2007ApJS..171..353S|uncertainty|   5.731   microns   | Broad-band measurement|03 27 04.4 -22 39 42.60 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
4|8.0 microns (IRAC)  | 89.9      |+/-9.9  | microJy            |3.81E+13|  8.99E-05|+/-9.90E-06|Jy|2007ApJS..171..353S|uncertainty|   7.872   microns   | Broad-band measurement|03 27 04.4 -22 39 42.60 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
5|5000 MHz            | 0.080     ||Jy                  |5.00E+09|  8.00E-02||Jy|1990PKS90.C...0000W|no uncertainty reported|    5000   MHz       | Broad-band measurement|03 24 51.5 -22 50 23 (B1950)| Integrated from scans|                                        |Homogenized from new and previously published data
6|4.85 GHz            | 131       |+/-13   |milliJy             |4.85E+09|  1.31E-01|+/-1.30E-02|Jy|1994ApJS...90..179G|rms noise|4.85       GHz       | Broad-band measurement|032702.3 -223956 (J2000)| Modelled datum|                                        |From new raw data; Corrected for contaminating sources
7|2700 MHz            | 0.200     ||Jy                  |2.70E+09|  2.00E-01||Jy|1990PKS90.C...0000W|no uncertainty reported|    2700   MHz       | Broad-band measurement|03 24 51.5 -22 50 23 (B1950)| Integrated from scans|                                        |Homogenized from new and previously published data
8|1.4GHz (VLA)        | 518.7     |+/-15.6 |milliJy             |1.40E+09|  5.19E-01|+/-1.56E-02|Jy|1998AJ....115.1693C|uncertainty|    1.40   GHz       | Broad-band measurement|03 27 4.46 -22 39 40.5 (J2000)| Flux integrated from map|                                        |From new raw data
9|408 MHz             | 1.98      |+/-0.10 |Jy                  |4.08E+08|  1.98E+00|+/-1.00E-01|Jy|1981MNRAS.194..693L|rms noise|408        MHz       | Broad-band measurement|032452.5 -225004 (B1950)| Modelled datum|                                        |From new raw data; Corrected for contaminating sources
10|408 MHz             | 1.980     ||Jy                  |4.08E+08|  1.98E+00||Jy|1990PKS90.C...0000W|no uncertainty reported|     408   MHz       | Broad-band measurement|03 24 51.5 -22 50 23 (B1950)| Integrated from scans|                                        |Homogenized from new and previously published data
11|365 MHz (Texas)     | 2.141     |+/-0.045|Jy                  |3.65E+08|  2.14E+00|+/-4.50E-02|Jy|1996AJ....111.1945D|internal error|365        MHz       | Broad-band measurement; obtained by interpolation over frequency|032452.633 -225003.63 (B1950)| Integrated from scans|Model:P;MFlag:+;EFlag:+;LFlag:+.        |From new raw data
12|74 MHz (VLA)        | 7.76      |+/-0.80 | Jy                 |7.38E+07|  7.76E+00|+/-8.00E-01|Jy|2007AJ....134.1245C|rms uncertainty|    73.8   MHz       | Broad-band measurement|03 27 04.13 -22 39 45.2 (J2000)| Flux integrated from map|Corrected for clean bias                |From new raw data
