
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-06-16T16:59:11PDT



Photometric Data for HS 1700+6416:[SSE2005] BX0561

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|U_n (WHT) AB        | 25.88     |+/-0.24 |mag                 |8.33E+14|  1.61E-07|+/-3.57E-08|Jy|2005ApJ...626..698S|estimated error|    0.36   microns   | Broad-band measurement|17 01 04.180 64 10 43.834 (J2000)| Flux integrated from map|                                        |From new raw data; derived from a flux in a different bandand a color
2|G (WHT) AB          | 24.84     |+/-0.18 |mag                 |6.38E+14|  4.21E-07|+/-6.93E-08|Jy|2005ApJ...626..698S|estimated error|    0.47   microns   | Broad-band measurement|17 01 04.180 64 10 43.834 (J2000)| Flux integrated from map|                                        |From new raw data; derived from a flux in a different bandand a color
3|G (WHT)             | 24.84     ||mag                 |6.38E+14|  4.21E-07||Jy|2006ApJ...647..128E|no uncertainty reported|    0.47   microns   | Broad-band measurement|| Flux in fixed aperture|                                        |Averaged from previously published data
4|H{alpha} (Keck II)  | 1.9E-17   |+/-0.6E-17|erg s^-1^ cm^-2^    |4.57E+14|  1.90E+06|+/-6.00E+05|Jy-Hz|2006ApJ...646..107E|uncertainty|    6563   A         | Line measurement; flux integrated over line; lines measured in emission|17 01 04.18 +64 10 43.83 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
5|R (WHT) AB          | 24.65     |+/-0.16 |mag                 |4.41E+14|  5.01E-07|+/-7.38E-08|Jy|2005ApJ...626..698S|estimated error|    0.68   microns   | Broad-band measurement|17 01 04.180 64 10 43.834 (J2000)| Flux integrated from map|                                        |From new raw data
6|J (Hale/WIRC)       | 22.30     ||mag                 |2.40E+14|  1.88E-06||Jy|2006ApJ...646..107E|no uncertainty reported|    1.25   microns   | Broad-band measurement|17 01 04.18 +64 10 43.83 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data; derived from aflux in a different band and a color
7|K_s (Hale/WIRC)     | 19.87     ||mag                 |1.39E+14|  7.55E-06||Jy|2006ApJ...646..107E|no uncertainty reported|    2.15   microns   | Broad-band measurement|17 01 04.18 +64 10 43.83 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data
8|K_s (P200) AB       | 21.84     |+/-0.19 |mag                 |1.39E+14|  6.67E-06|+/-1.19E-06|Jy|2005ApJ...626..698S|estimated error|    2.15   microns   | Broad-band measurement|17 01 04.180 64 10 43.834 (J2000)| Flux integrated from map|                                        |From new raw data; derived from a flux in a different bandand a color
9|3.6 microns IRAC AB | 21.54     |+/-0.10 |mag                 |8.33E+13|  8.79E-06|+/-8.09E-07|Jy|2005ApJ...626..698S|estimated error|     3.6   microns   | Broad-band measurement|17 01 04.180 64 10 43.834 (J2000)| Flux integrated from map|                                        |From new raw data
10|4.5 microns IRAC AB | 21.35     |+/-0.10 |mag                 |6.66E+13|  1.05E-05|+/-9.64E-07|Jy|2005ApJ...626..698S|estimated error|     4.5   microns   | Broad-band measurement|17 01 04.180 64 10 43.834 (J2000)| Flux integrated from map|                                        |From new raw data
11|5.8 microns IRAC AB | 21.19     |+/-0.10 |mag                 |5.17E+13|  1.21E-05|+/-1.12E-06|Jy|2005ApJ...626..698S|estimated error|     5.8   microns   | Broad-band measurement|17 01 04.180 64 10 43.834 (J2000)| Flux integrated from map|                                        |From new raw data
12|8.0 microns IRAC AB | 20.85     |+/-0.10 |mag                 |3.75E+13|  1.66E-05|+/-1.53E-06|Jy|2005ApJ...626..698S|estimated error|     8.0   microns   | Broad-band measurement|17 01 04.180 64 10 43.834 (J2000)| Flux integrated from map|                                        |From new raw data
