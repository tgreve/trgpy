

Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.


queryDateTime:2009-11-03T15:07:35PST






Photometric Data for MIPS8342 (z=1.5619)

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
4|R (KPNO)            | 1.171     ||microJy             |4.66E+14|  1.17E-06||Jy|2007ApJ...658..778Y|no uncertainty reported|    6440   A         | Broad-band measurement|171411.55 +601109.3 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data
5|R (Cousins) m_aper  | 23.84     |+/-0.08 |mag                 |4.65E+14|  8.91E-07|+/-6.56E-08|Jy|2004AJ....128....1F|based on count statistics only|6440       A         | Broad-band measurement|171411.471 +601109.31 (J2000)| Flux in fixed aperture|3-arcsecond aperture                    |From new raw data
6|R (Cousins) m_tot   | 23.50     |+/-0.12 |mag                 |4.65E+14|  1.22E-06|+/-1.35E-07|Jy|2004AJ....128....1F|based on count statistics only|6440       A         | Broad-band measurement|171411.471 +601109.31 (J2000)| Total flux|                                        |From new raw data
7|F160W (HST NICMOS)         | 20.26     ||mag                 |1.87E+14|  8.21E-06||Jy|2011ApJ...730..125Z|no uncertainty reported|      1.60 microns   | Broad-band measurement|| Flux integrated from map|                                        |From new raw data
8|F160W (HST NICMOS)         | 21.54     || mag                |1.86E+14|  2.53E-06||Jy|2008ApJ...680..232D|no uncertainty reported|      1.61 microns   | Broad-band measurement|17 14 11.45 +60 11 09.20 (J2000)| Flux integrated from map|                                        |From new raw data
9|3.6 microns (IRAC)  | 39        |+/-6    | microJy            |8.44E+13|  3.90E-05|+/-6.00E-06|Jy|2007ApJ...664..713S|uncertainty|   3.550   microns   | Broad-band measurement|| Flux in fixed aperture|7.3" diameter aperture                  |From reprocessed raw data
10|3.6 microns (IRAC)  | 38.01     |+/-4.54 |microJy             |8.42E+13|  3.80E-05|+/-4.54E-06|Jy|2005ApJS..161...41L|uncertainty|3.56       microns   | Broad-band measurement|171411.45 +601109.2 (J2000)| Flux in fixed aperture|Aperture =       4.92 arcsec.           |From new raw data
11|4.5 microns (IRAC)  | 57        |+/-4    | microJy            |6.67E+13|  5.70E-05|+/-4.00E-06|Jy|2007ApJ...664..713S|uncertainty|   4.493   microns   | Broad-band measurement|| Flux in fixed aperture|7.3" diameter aperture                  |From reprocessed raw data
12|4.5 microns (IRAC)  | 59.13     |+/-7.39 |microJy             |6.63E+13|  5.91E-05|+/-7.39E-06|Jy|2005ApJS..161...41L|uncertainty|4.52       microns   | Broad-band measurement|171411.45 +601109.2 (J2000)| Flux in fixed aperture|Aperture =       4.92 arcsec.           |From new raw data
13|5.8 microns (IRAC)  | 53        |+/-12   | microJy            |5.23E+13|  5.30E-05|+/-1.20E-05|Jy|2007ApJ...664..713S|uncertainty|   5.731   microns   | Broad-band measurement|| Flux in fixed aperture|7.3" diameter aperture                  |From reprocessed raw data
14|5.8 microns (IRAC)  ||<100.00    |microJy             |5.23E+13||1.00E-04|Jy|2005ApJS..161...41L|3sigma plate limit|5.73       microns   | Broad-band measurement|171411.45 +601109.2 (J2000)| Flux in fixed aperture|Aperture =       4.92 arcsec.           |From new raw data
17|8.0 microns (IRAC)  | 117.992   ||microJy             |3.81E+13|  1.18E-04||Jy|2007ApJ...658..778Y|no uncertainty reported|   7.872   microns   | Broad-band measurement|171411.55 +601109.3 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data
18|8.0 microns (IRAC)  | 119       |+/-19   | microJy            |3.81E+13|  1.19E-04|+/-1.90E-05|Jy|2007ApJ...664..713S|uncertainty|   7.872   microns   | Broad-band measurement|| Flux in fixed aperture|7.3" diameter aperture                  |From reprocessed raw data
19|8.0 microns (IRAC)  | 135.88    |+/-19.99|microJy             |3.79E+13|  1.36E-04|+/-2.00E-05|Jy|2005ApJS..161...41L|uncertainty|7.91       microns   | Broad-band measurement|171411.45 +601109.2 (J2000)| Flux in fixed aperture|Aperture =       4.92 arcsec.           |From new raw data
21|24 microns (MIPS)   | 1112.190  ||microJy             |1.27E+13|  1.11E-03||Jy|2007ApJ...658..778Y|no uncertainty reported|   23.68   microns   | Broad-band measurement|171411.55 +601109.3 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data; measurementmodified from published value
1|MIPS 24um           | 1.17     |+/-30%  |milliJy             |1.27E+13|  1.17E-03|+/-0.35E-03 |Jy|1996AJ....111.1431B|uncertainty|1.49       GHz       | Broad-band measurement| | Peak flux|                                        |From new raw data
2|MIPS 70um           | 10.7     |+/-1.4  |milliJy             |4.20E+12|  10.7E-03|+/-1.4E-03|Jy|2010Natur.464..733S|uncertainty|     71.42 microns   | Broad-band measurement|21 35 11.6 -01 02 52.0 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
23|70 microns (MIPS)   | 10.3      |+/-1.8  | milliJy            |4.20E+12|  1.03E-02|+/-1.80E-03|Jy|2007ApJ...664..713S|estimated error|   71.42   microns   | Broad-band measurement|| Flux in fixed aperture|3 pixel radius aperture                 |From reprocessed raw data
3|MIPS 160um          | 29.0     |+/-11.0 |milliJy             |1.92E+12|  29.0E-03|+/-11.0E-03|Jy|2009A&A...502..541E|3 sigma|     155.9 microns   | Broad-band measurement| | Flux in fixed aperture|                                        |From reprocessed raw data
4|MAMBO 1200um        | 0.98     |+/-0.52 |milliJy             |2.50E+11|  0.98E-03|+/-0.52E-03|Jy|2004MNRAS.354..779G|uncertainty|      1200 microns   | Broad-band measurement|16 37 06.7 +40 53 15 (J2000)| Flux integrated from map|S/N = 3.81                              |From new raw data
5|VLA 1.4GHz          | 0.18     |+/-0.03 |milliJy             |1.4E9   |  0.18E-03|+/-0.03E-03 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
6|GMRT 610MHz         | 0.86     |+/-0.11 |milliJy             |610.E6  |  0.86E-03|+/-0.11E-03 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
