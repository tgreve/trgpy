
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-12-16T05:10:18PST



Photometric Data for [HB89] 1413+117

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|0.5-8 keV (Chandra) | 3.3E-14   |+/-0.5E-14|ergs/cm^2^/s        |1.03E+18|  3.20E-09|+/-4.85E-10|Jy|2007ApJ...661...19P|uncertainty|    4.25   keV       | Broad-band measurement|| From fitting to map|Unabsorbed flux                         |From reprocessed raw data; NED frequency assigned tomid-point of band in keV
2|0.5-8 keV (Chandra) | 2.7E-14   |+/-0.7E-14|ergs/cm^2^/s        |1.03E+18|  2.62E-09|+/-6.80E-10|Jy|2007ApJ...661...19P|uncertainty|    4.25   keV       | Broad-band measurement|| From fitting to map|Unabsorbed flux                         |From reprocessed raw data; NED frequency assigned tomid-point of band in keV
3|0.5-8 keV (Chandra) | 0.90E-13  |+/-0.24E-13|erg/cm^2^/s         |1.03E+18|  8.74E-09|+/-2.33E-09|Jy|2012ApJ...744..111P|uncertainty|      4.25 keV       | Broad-band measurement|| Total flux|                                        |From reprocessed raw data; Extinction-corrected for MilkyWay; NED frequency assigned to mid-point of band in keV
4|0.4-8 keV (Chandra) | 1.0E-13   ||ergs/cm^2^/s        |1.02E+18|  9.80E-09||Jy|2004ApJ...605...45D|no uncertainty reported|    4.20   keV       | Broad-band measurement|| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
5|0.5-4.5 keV (XMM)   | -13.74    ||log(erg/cm^2^/s)    |6.05E+17|  3.01E-09||Jy|2011A&A...536A..84V|no uncertainty reported|      2.50 keV       | Broad-band measurement|14 15 46.2 +11 29 43 (J2000)| Flux integrated from map|                                        |Averaged from previously published data; NED frequencyassigned to mid-point of band in keV
6|FUV (GALEX) AB      ||>23.0841   |mag                 |1.95E+15||2.12E-06|Jy|2012GMSC..C...0000S|3 sigma|1538.6     A         | Broad-band measurement|213.94238407629 11.495397479235 (J2000)| Flux integrated from map|upper limit inside NUV Kron aperture    |From new raw data
7|FUV (GALEX) AB      | 25.1047   |+/-0.790978|mag                 |1.95E+15|  3.30E-07|+/-2.40E-07|Jy|2012GMSC..C...0000S|uncertainty|1538.6     A         | Broad-band measurement|213.94238407629 11.495397479235 (J2000)| Flux in fixed aperture|Flux in 7.5 arcsec diameter aperture    |From new raw data
8|1700 A (SDSS)       | -14.656   ||log(erg/cm^2^/s/A)  |1.76E+15|  2.13E-04||Jy|2011MNRAS.410..860A|no uncertainty reported|      1700 A         | Broad-band measurement|213.942673 +11.495402 (J2000)| Flux integrated from map|                                        |From reprocessed raw data
9|NUV (GALEX) AB      | 22.7936   |+/-0.261851|mag                 |1.29E+15|  2.77E-06|+/-6.68E-07|Jy|2012GMSC..C...0000S|uncertainty|2315.7     A         | Broad-band measurement|213.94238407629 11.495397479235 (J2000)| Flux integrated from map|Kron flux in elliptical aperture        |From new raw data
10|NUV (GALEX) AB      | 23.8775   |+/-0.309206|mag                 |1.29E+15|  1.02E-06|+/-2.91E-07|Jy|2012GMSC..C...0000S|uncertainty|2315.7     A         | Broad-band measurement|213.94238407629 11.495397479235 (J2000)| Flux in fixed aperture|Flux in 7.5 arcsec diameter aperture    |From new raw data
11|I (HST)             | 16.44     ||mag                 |3.68E+14|  6.40E-04||Jy|2011ApJ...738...96M|no uncertainty reported|     0.814 microns   | Broad-band measurement|| Not reported in paper|                                        |From reprocessed raw data
12|Y (UKIDSS)          | 15.74     |+/-0.15 |mag                 |2.91E+14|  1.04E-03|+/-1.44E-04|Jy|2010MNRAS.406.1583W|uncertainty|      1.03 microns   | Broad-band measurement|213.942670 +11.495402 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
13|J (UKIDSS)          | 15.37     |+/-0.15 |mag                 |2.40E+14|  1.11E-03|+/-1.53E-04|Jy|2010MNRAS.406.1583W|uncertainty|      1.25 microns   | Broad-band measurement|213.942670 +11.495402 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
14|F160W (HST/NICMOS)  | 20.527    |+/-0.037| mag                |1.87E+14|  6.69E-06|+/-2.28E-07|Jy|2007A&A...470..467C|internal error|       1.6 microns   | Broad-band measurement|| From fitting to map|                                        |From new raw data
15|F160W (HST/NIC2)    | 20.47     |+/-0.3  |mag                 |1.87E+14|  7.03E-06|+/-4.31E-06|Jy|2006ApJ...649..616P|typical accuracy|   1.606   microns   | Broad-band measurement|14 15 46.40 +11 29 41.4 (J2000)| From fitting to map|Host mag; extinction = 0.01             |From new raw data; Extinction-corrected for Milky Way
16|F160W (HST)         | 18.05     ||mag                 |1.87E+14|  6.29E-05||Jy|2011ApJ...742...93A|no uncertainty reported|      1.60 microns   | Broad-band measurement|| Not reported in paper|Unmagnified quasar mag                  |Averaged from previously published data
17|F160W (HST/NIC2)    | 18.41     ||mag                 |1.87E+14|  4.68E-05||Jy|2006ApJ...649..616P|no uncertainty reported|   1.606   microns   | Broad-band measurement|14 15 46.40 +11 29 41.4 (J2000)| From fitting to map|Quasar mag; extinction = 0.01           |From new raw data; Extinction-corrected for Milky Way
18|H (UKIDSS)          | 14.75     |+/-0.15 |mag                 |1.84E+14|  1.31E-03|+/-1.81E-04|Jy|2010MNRAS.406.1583W|uncertainty|      1.63 microns   | Broad-band measurement|213.942670 +11.495402 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
19|F180M (HST/NICMOS)  | 22.182    |+/-0.101| mag                |1.67E+14|  1.21E-06|+/-1.13E-07|Jy|2007A&A...470..467C|internal error|     1.795 microns   | Broad-band measurement|| From fitting to map|                                        |From new raw data
20|K (UKIDSS)          | 13.95     |+/-0.15 |mag                 |1.36E+14|  1.70E-03|+/-2.34E-04|Jy|2010MNRAS.406.1583W|uncertainty|      2.20 microns   | Broad-band measurement|213.942670 +11.495402 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
21|3.4 microns (WISE)  | 12.994    |+/-0.024|mag                 |8.82E+13|  1.96E-03|+/-4.34E-05|Jy|2012AJ....144...49W|uncertainty|       3.4 microns   | Broad-band measurement|213.942657 +11.495400 (J2000)| Not reported in paper|                                        |Averaged from previously published data
22|4.6 microns (WISE)  | 11.646    |+/-0.025|mag                 |6.52E+13|  3.77E-03|+/-8.69E-05|Jy|2012AJ....144...49W|uncertainty|       4.6 microns   | Broad-band measurement|213.942657 +11.495400 (J2000)| Not reported in paper|                                        |Averaged from previously published data
23|6.2 microns (IRS)   | 1.5E-21   ||W/cm^2^             |4.84E+13|  1.50E+09||Jy-Hz|2007ApJ...661L..25L|no uncertainty reported|     6.2   microns   | Line measurement; flux integrated over line; lines measured in emission|14 15 46.27 +11 29 43.40 (J2000)| Flux integrated from map|                                        |From new raw data
24|7.7 microns (IRS)   | 6.1E-21   ||W/cm^2^             |3.89E+13|  6.10E+09||Jy-Hz|2007ApJ...661L..25L|no uncertainty reported|     7.7   microns   | Line measurement; flux integrated over line; lines measured in emission|14 15 46.27 +11 29 43.40 (J2000)| Flux integrated from map|                                        |From new raw data
3|IRAS 12 microns     | |<93        |milliJy             |2.50E+13| |93.0E-03|Jy|1999ApJ...519..610D|3sisgma uncertainty reported| 12        microns   | Broad-band measurement|164502.36 +462625.5 (J2000)| Integrated from scans|                                        |Averaged from previously published data
25|12 microns (WISE)   | 7.747     |+/-0.020|mag                 |2.50E+13|  2.52E-02|+/-4.65E-04|Jy|2012AJ....144...49W|uncertainty|        12 microns   | Broad-band measurement|213.942657 +11.495400 (J2000)| Not reported in paper|                                        |Averaged from previously published data
26|22 microns (WISE)   | 5.404     |+/-0.030|mag                 |1.36E+13|  5.76E-02|+/-1.59E-03|Jy|2012AJ....144...49W|uncertainty|        22 microns   | Broad-band measurement|213.942657 +11.495400 (J2000)| Not reported in paper|                                        |Averaged from previously published data
6|IRAS 25 microns     | |<126.     |milliJy             |1.20E+13| |126.0E-03|Jy|1999ApJ...519..610D|3sigma uncertainty reported| 25        microns   | Broad-band measurement|164502.36 +462625.5 (J2000)| Integrated from scans|                                        |Averaged from previously published data
14|60 microns (IRAS)   | 230.0     |+/-38.0 |mJy                 |5.00E+12|230.0E-3|38.0E-03|Jy|2008A&A...477...55H|3rms uncertainty|     23.68 microns   | Broad-band measurement|14 00 57.530 +02 52 49.34 (J2000)| Flux in fixed aperture|6" radius aperture                      |From reprocessed raw data
15|100 microns (IRAS)  | 370.      |+/-78.  |mJy                 |3.00E+12|370.E-03|+/-78.E-03|Jy|1999ApJ...519..610D|3rms uncertainty| 20        cm        | Broad-band measurement|164502.36 +462625.5 (J2000)| Not reported in paper|                                        |Averaged from previously published data
27|[N II] 122 (CSO)    | 3.03E-18  |+/-0.29E-18|W/m^2^              |2.46E+12|  3.03E+08|+/-2.90E+07|Jy-Hz|2011ApJ...740L..29F|statistical error|       122 microns   | Line measurement; flux integrated over line; lines measured in emission|14 15 46.3 -11 29 44 (J2000)| Flux integrated from map|                                        |From new raw data
28|[N II] (IRAM)       ||<26.7      | Jy km/s            |1.46E+12||3.66E+07|Jy-Hz|2009ApJ...691L...1W|3 sigma|  1461.132 GHz       | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|                                        |From new raw data
29|CO (9-8) (CSO)      | 41.8      |+/-5.8  |Jy km/s             |1.04E+12|  4.07E+07|+/-5.64E+06|Jy-Hz|2009ApJ...705..112B|statistical error|   1036.91 GHz       | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|                                        |From new raw data
30|CO (8-7) (CSO)      | 51.4      |+/-4.7  |Jy km/s             |9.22E+11|  4.44E+07|+/-4.06E+06|Jy-Hz|2009ApJ...705..112B|statistical error|    921.80 GHz       | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|                                        |From new raw data
12|350 microns (SCUBA) | 189.0     |+/-56.0 |milliJy             |8.573E+11|189.0E-03|+/-56.0E-03|Jy|2007MNRAS.376.1073Z|3sigma uncertainty|     450   microns   | Broad-band measurement|02 39 51.9 -01 35 55 (J2000)| Flux integrated from map|                                        |From reprocessed raw data
31|350 microns (SHARC) | 0.293     |+/-0.014|Jy                  |8.57E+11|  2.93E-01|+/-1.40E-02|Jy|1999CIT...T00R....B|1 sigma|350        microns   | Broad-band measurement|141320.1 +114338. (B1950)| Flux integrated from map|                                        |From new raw data; OBJ_NAME modified from published value
32|[C I] (2-1) (CSO)   | 8.5       |+/-7.4  |Jy km/s             |8.09E+11|  6.45E+06|+/-5.62E+06|Jy-Hz|2009ApJ...705..112B|statistical error|    809.34 GHz       | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|                                        |From new raw data
33|CO (7-6) (CSO)      | 45.3      |+/-6.3  |Jy km/s             |8.07E+11|  3.43E+07|+/-4.77E+06|Jy-Hz|2009ApJ...705..112B|statistical error|    806.65 GHz       | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|                                        |From new raw data
34|CO (6-5) (CSO)      | 37.0      |+/-8.1  |Jy km/s             |6.91E+11|  2.40E+07|+/-5.25E+06|Jy-Hz|2009ApJ...705..112B|statistical error|    691.47 GHz       | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|                                        |From new raw data
16|450 microns (SCUBA) | 224.      |+/-38.  |milliJy             |6.66E+11|  224.E-03|+/-38.00E-03|Jy|2007MNRAS.376.1073Z|uncertainty|     450   microns   | Broad-band measurement|14 01 04.7 +02 52 28 (J2000)| Flux integrated from map|                                        |From reprocessed raw data
16|750 microns (SCUBA) | 44.0      |+/-8.0 |milliJy             |3.99E+11|  44.0E-03|+/-8.0E-03 |Jy|2007MNRAS.376.1073Z|no uncertainty reported|     850   microns   | Broad-band measurement|02 39 51.9 -01 35 55 (J2000)| Flux integrated from map|S/N = 19.9                              |From reprocessed raw data
35|HCO+(J=4-3) (PdBI)  | 0.54      |+/-0.09 |Jy km/s             |3.57E+11|  1.81E+05|+/-3.01E+04|Jy-Hz|2011ApJ...726...50R|uncertainty|  356.734  GHz       | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|                                        |From new raw data
36|^12CO (J=3-2) IRAM  | 30000     |+/-1700 |microJy             |3.46E+11|  3.00E-02|+/-1.70E-03|Jy|2006ApJ...645L..13R|uncertainty|345.7960   GHz       | Line measurement; flux integrated over line; lines measured in emission|| Peak flux|From 2003A&A...409L..41W                |Averaged from previously published data
37|CN(N=3-2) (PdBI)    | 1.94      |+/-0.24 | milliJy            |3.40E+11|  1.94E-03|+/-2.40E-04|Jy|2007ApJ...666..778R|uncertainty| 339.447   GHz       | Line measurement; flux integrated over line; lines measured in emission|| Peak flux|                                        |From new raw data
38|CN(N=3-2) (PdBI)    | 1.37      |+/-0.17 | Jy km/s            |3.40E+11|  5.11E+05|+/-6.34E+04|Jy-Hz|2007ApJ...666..778R|uncertainty| 2.55784             | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|                                        |From new raw data
39|^13^CO(3-2) (IRAM)  | 0.3       |+/-0.1  |Jy km/s             |3.31E+11|  1.49E+07|+/-4.97E+06|Jy-Hz|2010A&A...516A.111H|uncertainty|    330.59 GHz       | Line measurement; flux integrated over line; lines measured in emission|14 15 46.28 +11 29 44.0 (J2000)| Flux integrated from map|6.1" x 5.4" beam                        |From new raw data
26|1200 microns (MAMBO)| 16.0      |+/-2.0  | milliJy            |2.50E+11|  16.0E-03|+/-2.00E-03|Jy|2004MNRAS.354..779G|uncertainty|      1200 microns   | Broad-band measurement|16 36 50.3 +40 57 36 (J2000)| Flux integrated from map|S/N = 4.42                              |From new raw data
21|SCUBA 1350 microns  |           |<30.0   |milliJy             |2.22E+11|          |30.0E-03|Jy|1999ApJ...519..610D|3sigma uncertainty| 1350      microns   | Broad-band measurement|164502.36 +462625.5 (J2000)| Flux integrated from map|                                        |From new raw data
40|CO(1-0) (GBT)       | 1.406     |+/-0.053|Jy km/s             |1.15E+11|  1.52E+05|+/-5.73E+03|Jy-Hz|2011ApJ...739L..32R|uncertainty|   115.271 GHz       | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|Measured with Zpectrometer backend      |From new raw data
41|CO(1-0) (EVLA)      | 1.378     |+/-0.250|Jy km/s             |1.15E+11|  1.49E+05|+/-2.70E+04|Jy-Hz|2011ApJ...739L..32R|uncertainty|   115.271 GHz       | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|                                        |From new raw data
42|CO(1-0) (GBT)       | 1.358     |+/-0.065|Jy km/s             |1.15E+11|  1.47E+05|+/-7.02E+03|Jy-Hz|2011ApJ...739L..32R|uncertainty|   115.271 GHz       | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|Measured with Spectrometer backend      |From new raw data
43|92.9 GHz (PDBI/IRAM)     | 0.3       |+/-0.1  |milliJy             |9.29E+10|  3.00E-04|+/-1.00E-04|Jy|2010A&A...516A.111H|uncertainty|      92.9 GHz       | Broad-band measurement|14 15 46.28 +11 29 44.0 (J2000)| Flux integrated from map|6.1" x 5.4" beam                        |From new raw data
44|HCO+ (J=1-0) (VLA)  | 193       |+/-28   |microJy             |8.92E+10|  1.93E-04|+/-2.80E-05|Jy|2006ApJ...645L..13R|uncertainty| 89.1885   GHz       | Line measurement; flux integrated over line; lines measured in emission|| Peak flux|                                        |From new raw data
45|HCN (J=1-0) (VLA)   | 240       |+/-40   |microJy             |8.86E+10|  2.40E-04|+/-4.00E-05|Jy|2006ApJ...645L..13R|uncertainty| 88.6304   GHz       | Line measurement; flux integrated over line; lines measured in emission|| Peak flux|From 2003Natur.426..636S                |Averaged from previously published data
46|14.9 GHz (VLA)      | 0.56      |+/-0.18 |milliJy             |1.49E+10|  5.60E-04|+/-1.80E-04|Jy|1996AJ....111.1431B|uncertainty|14.9       GHz       | Broad-band measurement|| Peak flux|                                        |From new raw data
47|8.48 GHz (VLA)      | 0.98      |+/-0.08 |milliJy             |8.48E+09|  9.80E-04|+/-8.00E-05|Jy|1996AJ....111.1431B|uncertainty|8.48       GHz       | Broad-band measurement|| Peak flux|                                        |From new raw data
48|4.89 GHz (VLA)      | 1.95      |+/-0.13 |milliJy             |4.89E+09|  1.95E-03|+/-1.30E-04|Jy|1996AJ....111.1431B|uncertainty|4.89       GHz       | Broad-band measurement|| Peak flux|                                        |From new raw data
49|1.49 GHz (VLA)      | 7.68      |+/-0.50 |milliJy             |1.49E+09|  7.68E-03|+/-5.00E-04|Jy|1996AJ....111.1431B|uncertainty|1.49       GHz       | Broad-band measurement|| Peak flux|                                        |From new raw data
50|1.4GHz (VLA)        | 8.2       |+/-0.6  |milliJy             |1.40E+09|  8.20E-03|+/-6.00E-04|Jy|1998AJ....115.1693C|uncertainty|    1.40   GHz       | Broad-band measurement|14 15 46.09 +11 29 43.6 (J2000)| Flux integrated from map|                                        |From new raw data
