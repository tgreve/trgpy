
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-07-10T09:26:15PDT



Photometric Data for LEDA 2822840

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|3.6 microns (IRAC)  | 108.0     |+/-11.0 | microJy            |8.44E+13|  1.08E-04|+/-1.10E-05|Jy|2007ApJS..171..353S|uncertainty|   3.550   microns   | Broad-band measurement|01 54 55.8 -20 40 26.30 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
2|4.5 microns (IRAC)  | 165.0     |+/-17.0 | microJy            |6.67E+13|  1.65E-04|+/-1.70E-05|Jy|2007ApJS..171..353S|uncertainty|   4.493   microns   | Broad-band measurement|01 54 55.8 -20 40 26.30 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
3|5.8 microns (IRAC)  | 215.0     |+/-22.0 | microJy            |5.23E+13|  2.15E-04|+/-2.20E-05|Jy|2007ApJS..171..353S|uncertainty|   5.731   microns   | Broad-band measurement|01 54 55.8 -20 40 26.30 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
4|8.0 microns (IRAC)  | 415.0     |+/-42.0 | microJy            |3.81E+13|  4.15E-04|+/-4.20E-05|Jy|2007ApJS..171..353S|uncertainty|   7.872   microns   | Broad-band measurement|01 54 55.8 -20 40 26.30 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
5|39.9 GHz (ATCA)     | 5.1       |+/-1.5  |milliJy             |3.99E+10|  5.10E-03|+/-1.50E-03|Jy|2011ApJ...734L..25E|uncertainty|      39.9 GHz       | Broad-band measurement|| Flux integrated from map|                                        |From new raw data
6|4.85 GHz            | 115       |+/-12   |milliJy             |4.85E+09|  1.15E-01|+/-1.20E-02|Jy|1994ApJS...90..179G|rms noise|4.85       GHz       | Broad-band measurement|015455.3 -204020 (J2000)| Modelled datum|                                        |From new raw data; Corrected for contaminating sources
7|1.4GHz              | 453.1     |+/-13.6 |milliJy             |1.40E+09|  4.53E-01|+/-1.36E-02|Jy|1998AJ....115.1693C|uncertainty|    1.40   GHz       | Broad-band measurement|01 54 55.73 -20 40 26.9 (J2000)| Flux integrated from map|                                        |From new raw data
8|408 MHz             | 1.55      |+/-0.05 |Jy                  |4.08E+08|  1.55E+00|+/-5.00E-02|Jy|1981MNRAS.194..693L|rms noise|408        MHz       | Broad-band measurement|015234.3 -205508 (B1950)| Modelled datum|                                        |From new raw data; Corrected for contaminating sources
9|365 MHz (Texas)     | 1.582     |+/-0.038|Jy                  |3.65E+08|  1.58E+00|+/-3.80E-02|Jy|1996AJ....111.1945D|internal error|365        MHz       | Broad-band measurement; obtained by interpolation over frequency|015234.099 -205507.76 (B1950)| Integrated from scans|Model:P;MFlag:+;EFlag:+;LFlag:+.        |From new raw data
10|74 MHz (VLA)        | 3.10      |+/-0.31 | Jy                 |7.38E+07|  3.10E+00|+/-3.10E-01|Jy|2007AJ....134.1245C|rms uncertainty|    73.8   MHz       | Broad-band measurement|01 54 55.72 -20 40 25.6 (J2000)| Flux integrated from map|Corrected for clean bias                |From new raw data
