
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-07-10T03:57:34PDT



Photometric Data for COSMOS_53

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
22|24 microns (MIPS)   | 0.36      |+/-0.01 |milliJy             |1.27E+13|  0.36E-03|+/-0.01E-03|Jy|2010ApJ...716..348B|no uncertainty reported|     23.68 microns   | Broad-band measurement|150.1583900 2.1396030 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
5|250 microns (SPIRE)| 26.      |+/-3.0 |mJy             |1.199e+12| 26.0E-03|+/-3.0e-03 |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
6|350 microns (SPIRE)| 22.      |+/-3.0  |mJy             |8.565e+11|22.0E-03 |+/-3.0e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
