
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-04-05T08:15:36PDT



Photometric Data for RGJ131236.01+424044.1 (z=2.243)

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|R (Subaru)          | 24.7      |+/-0.3  |mag                 |4.76E+14|  4.11E-07|+/-1.14E-07|Jy|2006ApJS..167..103F|rms uncertainty|    6300   A         | Broad-band measurement|| Flux in fixed aperture|3" radius aperture                      |From new raw data
3|I (Cousins)         | 23.75     |+/-0.11 |mag                 |3.79E+14|  8.06E-07|+/-8.60E-08|Jy|2004ApJ...616...71S|1 sigma|    7900   A         | Broad-band measurement|| Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
4|z (Subaru)          | 24.3      |+/-0.5  |mag                 |3.26E+14|  4.17E-07|+/-1.92E-07|Jy|2006ApJS..167..103F|rms uncertainty|    9200   A         | Broad-band measurement|| Flux in fixed aperture|3" radius aperture                      |From new raw data
5|J (2MASS)           | 22.40     |+/-0.30 |mag                 |2.40E+14|  1.75E-06|+/-5.56E-07|Jy|2004ApJ...616...71S|1 sigma|    1.25   microns   | Broad-band measurement|| Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
6|K_s (2MASS)         | 20.50     |+/-0.27 |mag                 |1.38E+14|  4.21E-06|+/-1.19E-06|Jy|2004ApJ...616...71S|1 sigma|    2.17   microns   | Broad-band measurement|| Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
3|850 microns (SCUBA) |           |<3.3    |mJy             |3.53E+11|  |3.3E-03|Jy|2005MNRAS.358..149P|3sigma uncertainty|     850   microns   | Broad-band measurement|12 37 11.7 +62 22 12 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
7|850 microns (SCUBA) | 0.4       |+/-1.1  | milliJy            |3.53E+11|0.4E-03|+/-1.10E-03|Jy|2004ApJ...614..671C|1 sigma|       850 microns   | Broad-band measurement|131236.05 +424044.1 (J2000)| Flux integrated from map|                                        |From new raw data
5|1.4 GHz (VLA)       | 43.9      |+/-7.1  | microJy        |1.40E+09| 43.9E-06|+/-7.1E-06|Jy|2006MNRAS.371..963B|1 sigma|       1.4 GHz       | Broad-band measurement|16 36 55.767 +40 59 09.97 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
8|1.4 GHz (VLA)       | 54        |+/-10   |microJy             |1.40E+09|  5.40E-05|+/-1.00E-05|Jy|2006ApJS..167..103F|uncertainty|     1.4   GHz       | Broad-band measurement|13 12 36.066 +42 40 44.17 (J2000)| Flux integrated from map|Corrected to the sky; see paper         |From new raw data
