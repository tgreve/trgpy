


Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.





Photometric Data, HDF850.1, z=5.183 

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|F775W (HST/ACS) AB  |       |>24.6 |mag |3.86E+14 | |5.25e-07|Jy|2006ApJ...653...53B|3rms uncertainty reported|    7764   A         | Broad-band measurement|12 36 18.39 +62 15 50.1 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data; derived from a flux in a differentband and a color
2|3.6 microns (IRAC)  |       |<19.5 |uJy |8.44E+13 | |19.5E-06   |Jy|2011ApJ...728L...4H|3rms uncertainty       | | | | |
3|4.5 microns (IRAC)  |       |<17.6 |uJy |6.67E+13 | |17.6E-06   |Jy|2011ApJ...728L...4H|3rms uncertainty       | | | | |
4|5.8 microns (IRAC)  |       |<13.4 |uJy |5.23E+13 | |13.4E-06   |Jy|2009AJ....137.3884R|3rms uncertainty       | | | | |
5|8.0 microns (IRAC)  |       |<16.2 |uJy |3.85E+13 | |16.2E-06  |Jy|2009ApJ...699.1610H|3rms uncertainty       | | | | |
6|24um (Spitzer)      |       |<26.1 |uJy | 1.25E13 | |26.1E-6 |Jy |2003MNRAS.343..293M|3rms uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
7|24um (Spitzer)      | 28.2  |+/-4.4|uJy | 1.25E13 | 28.2E-6  |+/-4.4E-6 |Jy |2003MNRAS.343..293M|3rms uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
8|70 microns (MIPS)   |       |<2.0  |mJy |4.20E+12| |2.0E-03|Jy|2008ApJ...675..262R|2sigma uncertainty reported|     71.42 microns   | Broad-band measurement|14 01 04.96 +02 52 24.8 (J2000)| Flux in fixed aperture|                                        |From new raw data
9|100 microns (PACS)  |       |<1.18 |mJy |2.998e+12| |1.18E-03 |Jy|Reference          |3rms uncertainty       | | | | |
10|160 microns (PACS)  |       |<2.42 |mJy |1.874e+12| |2.42E-03 |Jy|Reference          |3rms uncertainty       | | | | |
11|250 microns (SPIRE) |       |<11.4 |mJy |1.199e+12| |11.4E-03 |Jy|Reference          |3rms uncertainty       | | | | |
12|350 microns (SPIRE) |       |<12.8 |mJy |8.57e+11 | |12.8E-03 |Jy|Reference          |3rms uncertainty       | | | | |
13|450 microns (SCUBA) |       |<21   |mJy |6.66E+11 | |21.0E-03 |Jy|2002MNRAS.331..495S|3rms uncertainty reported|     450   microns   | Broad-band measurement|140105.0 +025225 (J2000)| Flux integrated from map|                                        |From new raw data
14|500 microns (SPIRE) |       |<14.0 |mJy |5.996e+11| |14.0E-03 |Jy|Reference          |3rms uncertainty       | | | | |
15|850um (SCUBA)       | 7.0   |+/-0.4|mJy | 3.529E11| 7.0E-03  |+/-0.4E-3 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
16|850um (SCUBA)       | 5.9   |+/-0.3|mJy | 3.529E11| 5.9E-03  |+/-0.3E-3 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
17|1.3 mm (PdBI)      | 2.2   |+/-0.3|mJy |2.31E+11 | 2.2E-03|+/-0.3E-03|Jy|2006ApJ...640..228T|uncertainty|     1.3   mm        | Broad-band measurement| | Flux integrated from map|                                        |From new raw data
18|1.35 mm (SCUBA)    | 2.1   |+/-0.5|mJy |2.22E+11 | 2.1E-03|+/-0.5E-03|Jy|2006ApJ...640..228T|uncertainty|     1.3   mm        | Broad-band measurement| | Flux integrated from map|                                        |From new raw data
19|3.55 cm (VLA)      | 7.5   |+/-2.2|uJy |8.44E+09 | 7.5E-06  |+/-2.2E-06|Jy|2010A&A...518L..35I|uncertainty|      3.55 cm        | Broad-band measurement| | Flux integrated from map|                                        |From new raw data
20|1.4GHz (VLA)       | 16.73 |+/-4.25|uJy| 1.4E9   | 16.73E-6|+/-4.25E-6 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
21|1.4GHz (VLA)       |       |<15.9|uJy| 1.4E9   | |15.9E-6 |Jy |2003MNRAS.343..293M|3rms uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
