
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-06-16T17:10:41PDT



Photometric Data for [HB89] 2343+125:BX0389

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|G (WHT)             | 25.13     ||mag                 |6.38E+14|  3.22E-07||Jy|2006ApJ...647..128E|no uncertainty reported|    0.47   microns   | Broad-band measurement|| Flux in fixed aperture|                                        |Averaged from previously published data
2|H{beta} (VLT)       | 0.37E-16  |+/-0.05E-16|erg/s/cm^2^         |6.17E+14|  3.70E+06|+/-5.00E+05|Jy-Hz|2009ApJ...699.1660L|uncertainty|      4861 A         | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|                                        |From new raw data
3|R (Hale)            | 24.85     || mag                |4.76E+14|  3.54E-07||Jy|2007ApJ...670...15R|no uncertainty reported|      6300 A         | Broad-band measurement|| Not reported in paper|                                        |Averaged new and previously published data
4|H{alpha} (Keck II)  | 12.0E-17  |+/-0.4E-17|erg s^-1^ cm^-2^    |4.57E+14|  1.20E+07|+/-4.00E+05|Jy-Hz|2006ApJ...646..107E|uncertainty|    6563   A         | Line measurement; flux integrated over line; lines measured in emission|23 46 28.90 +12 47 33.55 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
5|H{alpha} (VLT)      | 21.0E-17  |+/-1.0E-17|erg/s/cm^2^         |4.57E+14|  2.10E+07|+/-1.00E+06|Jy-Hz|2009ApJ...706.1364F|uncertainty|      6563 A         | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|                                        |From new raw data
6|[S II] 6716 (VLT)   | 5.9E-16   |+/-0.1E-16|erg/s/cm^2^         |4.46E+14|  5.90E+07|+/-1.00E+06|Jy-Hz|2009ApJ...699.1660L|uncertainty|      6716 A         | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|                                        |From new raw data
7|[S II] 6731 (VLT)   | 7.5E-16   |+/-0.1E-16|erg/s/cm^2^         |4.45E+14|  7.50E+07|+/-1.00E+06|Jy-Hz|2009ApJ...699.1660L|uncertainty|      6731 A         | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|                                        |From new raw data
8|J (Hale/WIRC)       | 22.92     ||mag                 |2.40E+14|  1.06E-06||Jy|2006ApJ...646..107E|no uncertainty reported|    1.25   microns   | Broad-band measurement|23 46 28.90 +12 47 33.55 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data; derived from aflux in a different band and a color
9|F160W (HST) AB      | 23.11     |+/-0.10 |mag                 |1.87E+14|  2.07E-06|+/-1.91E-07|Jy|2011ApJ...731...65F|uncertainty|     1.603 microns   | Broad-band measurement|| Flux in fixed aperture|                                        |From new raw data
10|K_s (Hale/WIRC)     | 20.18     ||mag                 |1.39E+14|  5.68E-06||Jy|2006ApJ...646..107E|no uncertainty reported|    2.15   microns   | Broad-band measurement|23 46 28.90 +12 47 33.55 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data
11|CO(3-2) (PdBI)      |           |+/-0.15 |Jy km/s             |3.46E+11||+/-5.46E+04|Jy-Hz|2010Natur.463..781T|1 sigma|   345.998 GHz       | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|                                        |From new raw data
12|CO(3-2) (PdBI)      ||<0.27      | Jy km/s            |3.46E+11||9.82E+04|Jy-Hz|2008ApJ...680..246T|2 sigma|   345.796 GHz       | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|                                        |From new raw data
