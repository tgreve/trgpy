
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-05-28T01:50:15PDT



Photometric Data for PJ120207.6, z=2.4417

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
26|22 microns (WISE)  | 6.2       |+/-0.8|mJy           |1.36E+13|6.2E-03|0.8E-03|Jy|2012AJ....144...49W|3sigma limit|        22 microns   | Broad-band measurement|213.942657 +11.495400 (J2000)| Not reported in paper|                                        |Averaged from previously published data
1|250 microns (SPIRE) | 618.0     |+/-62.  |mJy         |1.199e+12|618.0E-03 |+/-62.0e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
1|250 microns (SPIRE) | 619.0     |+/-6.  |mJy         |1.199e+12|619.0E-03 |+/-6.0e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
3|350 microns (SPIRE) | 646.0     |+/-65.  |mJy         |8.565e+11|646.0E-03 |+/-65.0e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
3|350 microns (SPIRE) | 664.0     |+/-8.  |mJy         |8.565e+11|664.0E-03 |+/-8.0e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
5|350 microns (PLANCK) | 401.0    |+/-225.  |mJy        |8.57e+11|401.0E-03 |+/-225.0e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
5|500 microns (SPIRE) | 451.0     |+/-45.  |mJy         |5.996e+11|451.0E-03 |+/-45.0e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
5|500 microns (SPIRE) | 474.0     |+/-6.  |mJy         |5.996e+11|474.0E-03 |+/-6.0e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
9|850 microns (SCUBA) | 123.0     |+/-14. |milliJy       |3.53E+11|  123.E-03|+/-14.E-03 |Jy|2002MNRAS.331..495S|no uncertainty reported|     850   microns   | Broad-band measurement|140105.0 +025225 (J2000)| Flux integrated from map|                                        |From new raw data
2|1.1mm (AzTEC)        | 68.7 |+/-7.0| mJy  | 2.73E11| 68.7E-3| 7.9E-3 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
5|GISMO(2000.0um)     |  7.0   |+/-1.0 |mJy          |150.000E+9|7.0E-03 |+/-1.0E-03|Jy|2010ApJ...709..210K|uncertainty|      870  microns   | Broad-band measurement|16 35 55.67 +66 12 59.51 (J2000)| Flux integrated from map|                                        |From new raw data
5|VLA K-band 23.2GHz    |  140   |+/-8 |mJy          |23.1991E+9|140.0E-06 |+/-8E-06|Jy|2010ApJ...709..210K|uncertainty|      870  microns   | Broad-band measurement|16 35 55.67 +66 12 59.51 (J2000)| Flux integrated from map|                                        |From new raw data
14|1.4GHz (VLA)        | 2.01    |+/-0.121 |uJy  | 1.4E9   | 2.01E-3|+/-0.121E-3 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
