
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-07-10T06:40:50PDT



Photometric Data for [HB89] 1246-057

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|2-10 keV (XMM)      | -13.47    ||log(erg/s/cm^2^)    |1.45E+18|  2.34E-09||Jy|2010A&A...515A...2S|no uncertainty reported|      6.00 keV       | Broad-band measurement|| Modelled datum|                                        |From reprocessed raw data; NED frequency assigned tomid-point of band in keV
2|0.3-10 keV (XMM)    | 0.04E-12  ||erg cm^-2^ s^-1^    |1.25E+18|  3.20E-09||Jy|2005MNRAS.364..195P|no uncertainty reported|    5.15   keV       | Broad-band measurement|12 49 13.8 -05 59 18.0 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
3|0.5-2 keV           | 3.39E-14  |+/-0.85E-14|erg cm^-2^ s^-1^    |3.02E+17|  1.12E-08|+/-2.81E-09|Jy|2005MNRAS.360..610S|uncertainty|    1.25   keV       | Broad-band measurement|12 49 13.85 -05 59 19.4 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data;Extinction-corrected for Milky Way; NED frequency assigned tomid-point of band in keV
4|0.5-2 keV (XMM)     | -13.85    ||log(erg/s/cm^2^)    |3.02E+17|  4.68E-09||Jy|2010A&A...515A...2S|no uncertainty reported|      1.25 keV       | Broad-band measurement|| Modelled datum|                                        |From reprocessed raw data; NED frequency assigned tomid-point of band in keV
5|V                   | 16.7      ||mag                 |5.42E+14|  7.60E-04||Jy|2006ApJ...636..610R|no uncertainty reported|    5530   A         | Broad-band measurement|| Not reported in paper|                                        |Averaged from previously published data; Standard JohnsonUBVRI filters assumed
6|F702W (HST/WFPC2)   | 22.21     |+/-0.02 |mag                 |4.37E+14|  3.84E-06|+/-7.07E-08|Jy|2007ApJ...662..909K|uncertainty|    6862   A         | Broad-band measurement|| Flux in fixed aperture|                                        |From reprocessed raw data
7|J (AAO)             | 15.20     ||mag                 |2.50E+14|  1.36E-03||Jy|1982MNRAS.199..943H|no uncertainty reported|   1.20    microns   | Broad-band measurement|| Flux in fixed aperture|                                        |From new raw data; derived from a flux in a different bandand a color
8|H (AAO)             | 14.43     ||mag                 |1.83E+14|  1.74E-03||Jy|1982MNRAS.199..943H|no uncertainty reported|   1.64    microns   | Broad-band measurement|| Flux in fixed aperture|                                        |From new raw data; derived from a flux in a different bandand a color
9|K (AAO)             | 13.71     ||mag                 |1.37E+14|  2.13E-03||Jy|1982MNRAS.199..943H|no uncertainty reported|   2.19    microns   | Broad-band measurement|| Flux in fixed aperture|                                        |From new raw data
10|450 microns (SCUBA) | 81        |+/-12   |milliJy             |6.66E+11|  8.10E-02|+/-1.20E-02|Jy|2005MNRAS.360..610S|uncertainty|     450   microns   | Broad-band measurement|12 49 13.85 -05 59 19.4 (J2000)| Flux integrated from map|                                        |From new raw data
11|850 microns (SCUBA) | 7.2       |+/-1.4  |milliJy             |3.53E+11|  7.20E-03|+/-1.40E-03|Jy|2005MNRAS.360..610S|uncertainty|     850   microns   | Broad-band measurement|12 49 13.85 -05 59 19.4 (J2000)| Flux integrated from map|Original refcode=2001Sci...294.2516P    |Averaged from previously published data
12|114GHz | 0.65       |+/-0.02  |milliJy             |114.0E+09|  0.65E-03|+/-0.02E-03|Jy|2005MNRAS.360..610S|uncertainty|     850   microns   | Broad-band measurement|12 49 13.85 -05 59 19.4 (J2000)| Flux integrated from map|Original refcode=2001Sci...294.2516P    |Averaged from previously published data
