
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-06-16T17:12:49PDT



Photometric Data for [HB89] 2345+000:BX0482

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|G (WHT)             | 23.54     ||mag                 |6.38E+14|  1.39E-06||Jy|2006ApJ...647..128E|no uncertainty reported|    0.47   microns   | Broad-band measurement|| Flux in fixed aperture|                                        |Averaged from previously published data
2|H{alpha} (Keck II)  | 11.2E-17  |+/-0.3E-17|erg s^-1^ cm^-2^    |4.57E+14|  1.12E+07|+/-3.00E+05|Jy-Hz|2006ApJ...646..107E|uncertainty|    6563   A         | Line measurement; flux integrated over line; lines measured in emission|23 48 12.97 +00 25 46.34 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
3|H{alpha} (VLT)      | 23.2E-17  |+/-1.2E-17|erg/s/cm^2^         |4.57E+14|  2.32E+07|+/-1.20E+06|Jy-Hz|2009ApJ...706.1364F|uncertainty|      6563 A         | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|                                        |From new raw data
4|[S II] 6716 (VLT)   | 2.4E-16   |+/-0.1E-16|erg/s/cm^2^         |4.46E+14|  2.40E+07|+/-1.00E+06|Jy-Hz|2009ApJ...699.1660L|uncertainty|      6716 A         | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|                                        |From new raw data
5|[S II] 6731 (VLT)   | 3.1E-16   |+/-0.1E-16|erg/s/cm^2^         |4.45E+14|  3.10E+07|+/-1.00E+06|Jy-Hz|2009ApJ...699.1660L|uncertainty|      6731 A         | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|                                        |From new raw data
6|F160W (HST) AB      | 22.34     |+/-0.07 |mag                 |1.87E+14|  4.21E-06|+/-2.71E-07|Jy|2011ApJ...731...65F|uncertainty|     1.603 microns   | Broad-band measurement|| Flux in fixed aperture|                                        |From new raw data
