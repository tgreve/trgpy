
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-06-16T17:04:38PDT



Photometric Data for HS 1700+6416:[SSE2005] MD0069

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|U_n (WHT) AB        | 26.72     |+/-0.38 |mag                 |8.33E+14|  7.45E-08|+/-2.59E-08|Jy|2005ApJ...626..698S|estimated error|    0.36   microns   | Broad-band measurement|17 00 47.610 64 09 44.78 (J2000)| Flux integrated from map|                                        |From new raw data; derived from a flux in a different bandand a color
2|G (WHT) AB          | 25.22     |+/-0.18 |mag                 |6.38E+14|  2.96E-07|+/-5.01E-08|Jy|2005ApJ...626..698S|estimated error|    0.47   microns   | Broad-band measurement|17 00 47.610 64 09 44.78 (J2000)| Flux integrated from map|                                        |From new raw data; derived from a flux in a different bandand a color
3|G (WHT)             | 25.22     ||mag                 |6.38E+14|  2.96E-07||Jy|2006ApJ...647..128E|no uncertainty reported|    0.47   microns   | Broad-band measurement|| Flux in fixed aperture|                                        |Averaged from previously published data
4|H{alpha} (Keck II)  | 8.2E-17   |+/-0.9E-17|erg s^-1^ cm^-2^    |4.57E+14|  8.20E+06|+/-9.00E+05|Jy-Hz|2006ApJ...646..107E|uncertainty|    6563   A         | Line measurement; flux integrated over line; lines measured in emission|17 00 47.62 +64 09 44.78 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
5|R (WHT) AB          | 24.85     |+/-0.16 |mag                 |4.41E+14|  4.17E-07|+/-6.14E-08|Jy|2005ApJ...626..698S|estimated error|    0.68   microns   | Broad-band measurement|17 00 47.610 64 09 44.78 (J2000)| Flux integrated from map|                                        |From new raw data
6|J (Hale/WIRC)       | 22.65     ||mag                 |2.40E+14|  1.36E-06||Jy|2006ApJ...646..107E|no uncertainty reported|    1.25   microns   | Broad-band measurement|17 00 47.62 +64 09 44.78 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data; derived from aflux in a different band and a color
7|K_s (Hale/WIRC)     | 20.05     ||mag                 |1.39E+14|  6.40E-06||Jy|2006ApJ...646..107E|no uncertainty reported|    2.15   microns   | Broad-band measurement|17 00 47.62 +64 09 44.78 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data
8|K_s (P200) AB       | 21.80     |+/-0.20 |mag                 |1.39E+14|  6.92E-06|+/-1.27E-06|Jy|2005ApJ...626..698S|estimated error|    2.15   microns   | Broad-band measurement|17 00 47.610 64 09 44.78 (J2000)| Flux integrated from map|                                        |From new raw data; derived from a flux in a different bandand a color
9|3.6 microns IRAC AB | 21.13     |+/-0.03 |mag                 |8.33E+13|  1.28E-05|+/-3.54E-07|Jy|2005ApJ...626..698S|estimated error|     3.6   microns   | Broad-band measurement|17 00 47.610 64 09 44.78 (J2000)| Flux integrated from map|                                        |From new raw data
10|4.5 microns IRAC AB | 20.89     |+/-0.04 |mag                 |6.66E+13|  1.60E-05|+/-5.89E-07|Jy|2005ApJ...626..698S|estimated error|     4.5   microns   | Broad-band measurement|17 00 47.610 64 09 44.78 (J2000)| Flux integrated from map|                                        |From new raw data
11|5.8 microns IRAC AB | 20.59     |+/-0.07 |mag                 |5.17E+13|  2.11E-05|+/-1.36E-06|Jy|2005ApJ...626..698S|estimated error|     5.8   microns   | Broad-band measurement|17 00 47.610 64 09 44.78 (J2000)| Flux integrated from map|                                        |From new raw data
12|8.0 microns IRAC AB | 20.63     |+/-0.11 |mag                 |3.75E+13|  2.03E-05|+/-2.06E-06|Jy|2005ApJ...626..698S|estimated error|     8.0   microns   | Broad-band measurement|17 00 47.610 64 09 44.78 (J2000)| Flux integrated from map|                                        |From new raw data
13|CO(3-2) (PdBI)      ||<0.06      |Jy km/s             |3.46E+11|  1.47E+05|2.10E+04|Jy-Hz|2010Natur.463..781T|3 sigma|   345.998 GHz       | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|                                        |From new raw data
