\queryDateTime = 2018-11-24T07:06:24PST
\source = /hydra/workarea/irsaviewer/temp_files/IpacTableFromSource1766008363458859407.tbl
\QUERY_STATUS = OK
\CatalogTargetColName = Coordinates Targeted
\Description = Published and Homogenized [Frequency, Flux Dens...
\LINK = http://ned.ipac.caltech.edu/cgi-bin/datasearch?sea
\
z=0.01813
|No.    |Observed Passband   |Photometry Measurement|Uncertainty  |Units             |Frequency |Flux Densit y|Upper limit of uncertainty |Lower limit of uncertainty|Upper limit of Flux Density  |Lower limit of Flux Density |NED Uncertainty |NED Units |Refcode              |Significance                  |Published frequency |Frequency Mode                                                                               |Coordinates Targeted              |Spatial Mode                                               |Qualifiers                                |Comments                                          
|int    |char                |double                |char         |char              |double    |double       |double                     |double                    |double                       |double                      |char            |char      |char                 |char                          |char                |char                                                                                         |char                              |char                                                       |char                                      |char                                              
|       |                    |                      |             |                  |Hz        |Jy           |                           |                          |                             |                            |                |          |                     |                              |                    |                                                                                             |                                  |                                                           |                                          |                                                  
|       |                    |                      |             |                  |          |             |                           |                          |                             |                            |                |          |                     |                              |                    |                                                                                             |                                  |                                                           |                                          |                                                  
 1      |2-10 keV (ASCA)     |1.1E-13               |             |ergs/s/cm^2^      |1.45E+18  |7.59E-09     |                           |                          |                             |                            |                | Jy       | 2001ApJS..133....1U |no uncertainty reported       | 6.00 keV           | Broad-band measurement                                                                      | 233.7458 +23.4932 (J2000)        |Flux integrated from map                                   |                                          |From reprocessed raw data; Extinction-corrected for MilkyWay; NED frequency assigned to mid-point of band in keV                                                    
 2      |2-10 keV (Suzaku)   |9.8E-14               |+/-0.24E-13  |erg/s/cm^2^       |1.45E+18  |6.76E-09     |1.66E-09                   |1.66E-09                  |                             |                            | +/-1.66E-09    | Jy       | 2009ApJ...691..261T |uncertainty                   | 6.00 keV           | Broad-band measurement                                                                      |                                  |Modelled datum                                             |                                          |From new raw data; NED frequency assigned to mid-point ofband in keV                                                                                                
 3      |2-10 keV            |1.1E-13               |+/-0.18E-13  |erg/s/cm^2^       |1.45E+18  |7.38E-09     |1.24E-09                   |1.24E-09                  |                             |                            | +/-1.24E-09    | Jy       | 2011ApJ...729...52L |uncertainty                   | 6.00 keV           | Broad-band measurement                                                                      |                                  |Modelled datum                                             |                                          |From reprocessed raw data; NED frequency assigned tomid-point of band in keV                                                                                        
 4      |2-7 keV (Chandra)   |6.6E-14               |             |erg/s/cm^2^       |1.09E+18  |6.06E-09     |                           |                          |                             |                            |                | Jy       | 2011A&A...529A.106I |no uncertainty reported       | 4.50 keV           | Broad-band measurement                                                                      |                                  |Modelled datum                                             |                                          |From reprocessed raw data; NED frequency assigned tomid-point of band in keV                                                                                        
 5      |0.7-7 keV (ASCA)    |2.1E-13               |             |ergs/s/cm^2^      |9.31E+17  |2.26E-08     |                           |                          |                             |                            |                | Jy       | 2001ApJS..133....1U |no uncertainty reported       | 3.85 keV           | Broad-band measurement                                                                      | 233.7458 +23.4932 (J2000)        |Flux integrated from map                                   |                                          |From reprocessed raw data; Extinction-corrected for MilkyWay; NED frequency assigned to mid-point of band in keV                                                    
 6      |EO IPC (0.1-4.5 keV)|4.6E+01               |             |nJy               |3.87E+17  |4.57E-08     |                           |                          |                             |                            |                | Jy       | 1996MNRAS.278.1049R |no uncertainty reported       | 1.6        keV     | Broad-band measurement; broad-band flux derived by integration over spectrum; synthetic band| 153457.22 +233011.40 (J2000)     |Integrated from scans                                      |                                          |Homogenized from previously published data                                                                                                                          
 7      |0.7-2 keV (ASCA)    |1.4E-13               |             |ergs/s/cm^2^      |3.26E+17  |4.29E-08     |                           |                          |                             |                            |                | Jy       | 2001ApJS..133....1U |no uncertainty reported       | 1.35 keV           | Broad-band measurement                                                                      | 233.7458 +23.4932 (J2000)        |Flux integrated from map                                   |                                          |From reprocessed raw data; Extinction-corrected for MilkyWay; NED frequency assigned to mid-point of band in keV                                                    
 8      |0.5-2 keV (Suzaku)  |6.6E-14               |+/-0.10E-13  |erg/s/cm^2^       |3.02E+17  |2.19E-08     |3.31E-09                   |3.31E-09                  |                             |                            | +/-3.31E-09    | Jy       | 2009ApJ...691..261T |uncertainty                   | 1.25 keV           | Broad-band measurement                                                                      |                                  |Modelled datum                                             |                                          |From new raw data; NED frequency assigned to mid-point ofband in keV                                                                                                
 9      |0.5-2 keV (Chandra) |2.7E-14               |             |erg/s/cm^2^       |3.02E+17  |8.94E-09     |                           |                          |                             |                            |                | Jy       | 2011A&A...529A.106I |no uncertainty reported       | 1.25 keV           | Broad-band measurement                                                                      |                                  |Modelled datum                                             |                                          |From reprocessed raw data; NED frequency assigned tomid-point of band in keV                                                                                        
 10     |FUV (GALEX) AB      |1.9E+01               |+/-0.12      |mag               |1.96E+15  |9.42E-05     |1.01E-05                   |1.01E-05                  |                             |                            | +/-1.01E-05    | Jy       | 2014ApJS..212...18B |uncertainty                   | 1531   A           | Broad-band measurement                                                                      | 233.73850000 23.50317000 (J2000) |Flux in fixed aperture                                     |  80"x36" aperture; PSF corr              |From new raw data                                                                                                                                                   
 11     |FUV (GALEX) AB      |1.9E+01               |+/-0.12      |mag               |1.96E+15  |1.36E-04     |1.45E-05                   |1.45E-05                  |                             |                            | +/-1.45E-05    | Jy       | 2014ApJS..212...18B |uncertainty                   | 1531   A           | Broad-band measurement                                                                      | 233.73850000 23.50317000 (J2000) |Flux in fixed aperture                                     |  80"x36" aperture; PSF corr              |From new raw data; Extinction-corrected for Milky Way                                                                                                               
 12     |UVW2 (Swift) AB     |1.8E+01               |+/-0.10      |mag               |1.48E+15  |2.38E-04     |2.19E-05                   |2.19E-05                  |                             |                            | +/-2.19E-05    | Jy       | 2014ApJS..212...18B |uncertainty                   | 2026   A           | Broad-band measurement                                                                      | 233.73850000 23.50317000 (J2000) |Flux in fixed aperture                                     |  80"x36" aperture                        |From new raw data                                                                                                                                                   
 13     |UVW2 (Swift) AB     |1.8E+01               |+/-0.10      |mag               |1.48E+15  |3.46E-04     |3.18E-05                   |3.18E-05                  |                             |                            | +/-3.18E-05    | Jy       | 2014ApJS..212...18B |uncertainty                   | 2026   A           | Broad-band measurement                                                                      | 233.73850000 23.50317000 (J2000) |Flux in fixed aperture                                     |  80"x36" aperture                        |From new raw data; Extinction-corrected for Milky Way                                                                                                               
 14     |NUV (GALEX) AB      |1.8E+01               |+/-0.10      |mag               |1.31E+15  |3.13E-04     |2.88E-05                   |2.88E-05                  |                             |                            | +/-2.88E-05    | Jy       | 2014ApJS..212...18B |uncertainty                   | 2286   A           | Broad-band measurement                                                                      | 233.73850000 23.50317000 (J2000) |Flux in fixed aperture                                     |  80"x36" aperture; PSF corr              |From new raw data                                                                                                                                                   
 15     |NUV (GALEX) AB      |1.7E+01               |+/-0.10      |mag               |1.31E+15  |4.53E-04     |4.17E-05                   |4.17E-05                  |                             |                            | +/-4.17E-05    | Jy       | 2014ApJS..212...18B |uncertainty                   | 2286   A           | Broad-band measurement                                                                      | 233.73850000 23.50317000 (J2000) |Flux in fixed aperture                                     |  80"x36" aperture; PSF corr              |From new raw data; Extinction-corrected for Milky Way                                                                                                               
 16     |u (SDSS) AB         |1.5E+01               |+/-0.05      |mag               |8.44E+14  |2.32E-03     |1.07E-04                   |1.07E-04                  |                             |                            | +/-1.07E-04    | Jy       | 2014ApJS..212...18B |uncertainty                   | 3551   A           | Broad-band measurement                                                                      | 233.73850000 23.50317000 (J2000) |Flux in fixed aperture                                     |  80"x36" aperture                        |From new raw data                                                                                                                                                   
 17     |u (SDSS) AB         |1.5E+01               |+/-0.05      |mag               |8.44E+14  |2.85E-03     |1.31E-04                   |1.31E-04                  |                             |                            | +/-1.31E-04    | Jy       | 2014ApJS..212...18B |uncertainty                   | 3551   A           | Broad-band measurement                                                                      | 233.73850000 23.50317000 (J2000) |Flux in fixed aperture                                     |  80"x36" aperture                        |From new raw data; Extinction-corrected for Milky Way                                                                                                               
 18     |U_T (VATT)          |1.4E+01               |+/-0.023     |mag               |8.19E+14  |3.32E-03     |6.98E-05                   |6.98E-05                  |                             |                            | +/-6.98E-05    | Jy       | 2005ApJ...630..784T |uncertainty                   | 3660   A           | Broad-band measurement                                                                      | 15 34 56.33 +23 29 33.8 (J2000)  |Total flux                                                 |                                          |From new raw data; derived from a flux in a different bandand a color; Standard Johnson UBVRI filters assumed                                                       
 19     |U (U_T)             |1.4E+01               |+/-0.15      |mag               |8.19E+14  |3.55E-03     |5.09E-04                   |5.09E-04                  |                             |                            | +/-5.09E-04    | Jy       | 1991RC3.9.C...0000d |rms uncertainty               | 3660       A       | Broad-band measurement                                                                      | 153247.3 +234006 (B1950)         |From multi-aperture data                                   |                                          |Homogenized from new and previously published data; StandardJohnson UBVRI filters assumed                                                                           
 20     |U (U_T^0)           |1.4E+01               |             |mag               |8.19E+14  |5.13E-03     |                           |                          |                             |                            |                | Jy       | 1991RC3.9.C...0000d |no uncertainty reported       | 3660       A       | Broad-band measurement                                                                      | 153247.3 +234006 (B1950)         |From multi-aperture data                                   |                                          |Homogenized from new and previously published data;Extinction-corrected for internal and Milky Way and K-correction applied; Standard Johnson UBVRI filters assumed 
 22     |103a-O (POSS-I O)   |1.4E+01               |             |mag               |7.40E+14  |6.44E-03     |                           |                          |                             |                            |                | Jy       | 2006ApJ...639...37K |no uncertainty reported       | 4050   A           | Broad-band measurement                                                                      | 153457.1 +233007 (J2000)         |Flux integrated from map                                   |                                          |Averaged new and previously published data                                                                                                                          
 25     |m_p                 |1.4E+01               |+/-0.4       |mag               |6.81E+14  |7.40E-03     |3.30E-03                   |3.30E-03                  |                             |                            | +/-3.30E-03    | Jy       | 1963CGCG2.C...0000Z |rms noise                     | 4400       A       | Broad-band measurement                                                                      | 153248.0 +234000. (B1950)        |Estimated by eye                                           |                                          |From new raw data                                                                                                                                                   
 26     |B_T (VATT)          |1.4E+01               |+/-0.011     |mag               |6.81E+14  |1.06E-02     |1.07E-04                   |1.07E-04                  |                             |                            | +/-1.07E-04    | Jy       | 2005ApJ...630..784T |uncertainty                   | 4400   A           | Broad-band measurement                                                                      | 15 34 56.33 +23 29 33.8 (J2000)  |Total flux                                                 |                                          |From new raw data; Standard Johnson UBVRI filters assumed                                                                                                           
 27     |B (UH)              |1.4E+01               |+/-0.07      |mag               |6.81E+14  |1.07E-02     |6.90E-04                   |6.90E-04                  |                             |                            | +/-6.90E-04    | Jy       | 2000ApJ...529..170S |uncertainty                   | 4400   A           | Broad-band measurement                                                                      | 15 34 57.3 +23 30 11.9 (J2000)   |Flux in fixed aperture                                     |                                          |From new raw data                                                                                                                                                   
 28     |B (UH)              |1.8E+01               |+/-0.1       |mag               |6.81E+14  |3.89E-04     |3.58E-05                   |3.58E-05                  |                             |                            | +/-3.58E-05    | Jy       | 2000ApJ...529..170S |uncertainty                   | 4400   A           | Broad-band measurement                                                                      | 15 34 57.3 +23 30 11.9 (J2000)   |Flux in fixed aperture                                     |  Nuclear mag                             |From new raw data                                                                                                                                                   
 29     |B (B_T)             |1.4E+01               |+/-0.14      |mag               |6.81E+14  |1.13E-02     |1.56E-03                   |1.56E-03                  |                             |                            | +/-1.56E-03    | Jy       | 1991RC3.9.C...0000d |rms uncertainty               | 4400       A       | Broad-band measurement                                                                      | 153247.3 +234006 (B1950)         |From multi-aperture data                                   |                                          |Homogenized from new and previously published data; StandardJohnson UBVRI filters assumed                                                                           
 30     |B (m_B)             |1.4E+01               |+/-0.20      |mag               |6.81E+14  |1.17E-02     |2.37E-03                   |2.37E-03                  |                             |                            | +/-2.37E-03    | Jy       | 1991RC3.9.C...0000d |rms uncertainty               | 4400       A       | Broad-band measurement                                                                      | 153247.3 +234006 (B1950)         |Multiple methods                                           |                                          |Homogenized from new and previously published data; StandardJohnson UBVRI filters assumed                                                                           
 31     |B (B_T^0)           |1.4E+01               |             |mag               |6.81E+14  |1.53E-02     |                           |                          |                             |                            |                | Jy       | 1991RC3.9.C...0000d |no uncertainty reported       | 4400       A       | Broad-band measurement                                                                      | 153247.3 +234006 (B1950)         |Multiple methods                                           |                                          |Homogenized from new and previously published data;Extinction-corrected for internal and Milky Way and K-correction applied; Standard Johnson UBVRI filters assumed 
 32     |g (SDSS) AB         |1.4E+01               |+/-0.05      |mag               |6.40E+14  |1.04E-02     |4.81E-04                   |4.81E-04                  |                             |                            | +/-4.81E-04    | Jy       | 2014ApJS..212...18B |uncertainty                   | 4681   A           | Broad-band measurement                                                                      | 233.73850000 23.50317000 (J2000) |Flux in fixed aperture                                     |  80"x36" aperture                        |From new raw data                                                                                                                                                   
 33     |g (SDSS) AB         |1.4E+01               |+/-0.05      |mag               |6.40E+14  |1.23E-02     |5.65E-04                   |5.65E-04                  |                             |                            | +/-5.65E-04    | Jy       | 2014ApJS..212...18B |uncertainty                   | 4681   A           | Broad-band measurement                                                                      | 233.73850000 23.50317000 (J2000) |Flux in fixed aperture                                     |  80"x36" aperture                        |From new raw data; Extinction-corrected for Milky Way                                                                                                               
 37     |V_T (VATT)          |1.3E+01               |+/-0.018     |mag               |5.42E+14  |1.93E-02     |3.17E-04                   |3.17E-04                  |                             |                            | +/-3.17E-04    | Jy       | 2005ApJ...630..784T |uncertainty                   | 5530   A           | Broad-band measurement                                                                      | 15 34 56.33 +23 29 33.8 (J2000)  |Total flux                                                 |                                          |From new raw data; derived from a flux in a different bandand a color; Standard Johnson UBVRI filters assumed                                                       
 38     |V (V_T)             |1.3E+01               |+/-0.14      |mag               |5.42E+14  |1.91E-02     |2.69E-03                   |2.69E-03                  |                             |                            | +/-2.69E-03    | Jy       | 1991RC3.9.C...0000d |rms uncertainty               | 5530       A       | Broad-band measurement                                                                      | 153247.3 +234006 (B1950)         |From multi-aperture data                                   |                                          |Homogenized from new and previously published data; StandardJohnson UBVRI filters assumed                                                                           
 39     |V (V_T^0)           |1.3E+01               |             |mag               |5.42E+14  |2.38E-02     |                           |                          |                             |                            |                | Jy       | 1991RC3.9.C...0000d |no uncertainty reported       | 5530       A       | Broad-band measurement                                                                      | 153247.3 +234006 (B1950)         |From multi-aperture data                                   |                                          |Homogenized from new and previously published data;Extinction-corrected for internal and Milky Way and K-correction applied; Standard Johnson UBVRI filters assumed 
 40     |r (SDSS) AB         |1.3E+01               |+/-0.05      |mag               |4.86E+14  |2.23E-02     |1.03E-03                   |1.03E-03                  |                             |                            | +/-1.03E-03    | Jy       | 2014ApJS..212...18B |uncertainty                   | 6165   A           | Broad-band measurement                                                                      | 233.73850000 23.50317000 (J2000) |Flux in fixed aperture                                     |  80"x36" aperture                        |From new raw data; Extinction-corrected for Milky Way                                                                                                               
 41     |r (SDSS) AB         |1.3E+01               |+/-0.05      |mag               |4.86E+14  |2.00E-02     |9.22E-04                   |9.22E-04                  |                             |                            | +/-9.22E-04    | Jy       | 2014ApJS..212...18B |uncertainty                   | 6165   A           | Broad-band measurement                                                                      | 233.73850000 23.50317000 (J2000) |Flux in fixed aperture                                     |  80"x36" aperture                        |From new raw data                                                                                                                                                   
 44     |H{alpha} (WHT)      |3.1E-14               |+/-15  %     |ergs/s/cm^2^/A    |4.57E+14  |4.46E-02     |6.69E-03                   |6.69E-03                  |                             |                            | +/-6.69E-03    | Jy       | 2004ApJ...602..181C |uncertainty                   | 6563   A           | Line measurement; flux integrated over line; lines measured in emission                     |                                  |Flux integrated from map                                   |  Circumnuclear flux                      |From new raw data                                                                                                                                                   
 48     |R_T (VATT)          |1.2E+01               |+/-0.020     |mag               |4.33E+14  |2.97E-02     |5.58E-04                   |5.58E-04                  |                             |                            | +/-5.58E-04    | Jy       | 2005ApJ...630..784T |uncertainty                   | 6930   A           | Broad-band measurement                                                                      | 15 34 56.33 +23 29 33.8 (J2000)  |Total flux                                                 |                                          |From new raw data; derived from a flux in a different bandand a color; Standard Johnson UBVRI filters assumed                                                       
 49     |i (SDSS) AB         |1.3E+01               |+/-0.05      |mag               |4.01E+14  |2.94E-02     |1.35E-03                   |1.35E-03                  |                             |                            | +/-1.35E-03    | Jy       | 2014ApJS..212...18B |uncertainty                   | 7480   A           | Broad-band measurement                                                                      | 233.73850000 23.50317000 (J2000) |Flux in fixed aperture                                     |  80"x36" aperture                        |From new raw data                                                                                                                                                   
 50     |i (SDSS) AB         |1.3E+01               |+/-0.05      |mag               |4.01E+14  |3.19E-02     |1.47E-03                   |1.47E-03                  |                             |                            | +/-1.47E-03    | Jy       | 2014ApJS..212...18B |uncertainty                   | 7480   A           | Broad-band measurement                                                                      | 233.73850000 23.50317000 (J2000) |Flux in fixed aperture                                     |  80"x36" aperture                        |From new raw data; Extinction-corrected for Milky Way                                                                                                               
 51     |I (UH)              |1.2E+01               |+/-0.07      |mag               |3.79E+14  |3.21E-02     |2.07E-03                   |2.07E-03                  |                             |                            | +/-2.07E-03    | Jy       | 2000ApJ...529..170S |uncertainty                   | 7900   A           | Broad-band measurement                                                                      | 15 34 57.3 +23 30 11.9 (J2000)   |Flux in fixed aperture                                     |                                          |From new raw data                                                                                                                                                   
 52     |I (UH)              |1.5E+01               |+/-0.1       |mag               |3.79E+14  |3.36E-03     |3.10E-04                   |3.10E-04                  |                             |                            | +/-3.10E-04    | Jy       | 2000ApJ...529..170S |uncertainty                   | 7900   A           | Broad-band measurement                                                                      | 15 34 57.3 +23 30 11.9 (J2000)   |Flux in fixed aperture                                     |  Nuclear mag                             |From new raw data                                                                                                                                                   
 53     |z (SDSS) AB         |1.2E+01               |+/-0.05      |mag               |3.36E+14  |3.95E-02     |1.82E-03                   |1.82E-03                  |                             |                            | +/-1.82E-03    | Jy       | 2014ApJS..212...18B |uncertainty                   | 8931   A           | Broad-band measurement                                                                      | 233.73850000 23.50317000 (J2000) |Flux in fixed aperture                                     |  80"x36" aperture                        |From new raw data; Extinction-corrected for Milky Way                                                                                                               
 54     |z (SDSS) AB         |1.2E+01               |+/-0.05      |mag               |3.36E+14  |3.71E-02     |1.71E-03                   |1.71E-03                  |                             |                            | +/-1.71E-03    | Jy       | 2014ApJS..212...18B |uncertainty                   | 8931   A           | Broad-band measurement                                                                      | 233.73850000 23.50317000 (J2000) |Flux in fixed aperture                                     |  80"x36" aperture                        |From new raw data                                                                                                                                                   
 55     |J (ESO/SPM)         |2.8E+01               |+/-1.85      |milliJy           |2.50E+14  |2.78E-02     |1.85E-03                   |1.85E-03                  |                             |                            | +/-1.85E-03    | Jy       | 1995ApJ...453..616S |rms uncertainty               | 1.198      microns | Broad-band measurement                                                                      | 153246.8 +234007 (B1950)         |Flux in fixed aperture                                     |  15" aperture                            |From new raw data                                                                                                                                                   
 56     |J (2MASS) AB        |1.2E+01               |+/-0.05      |mag               |2.43E+14  |6.12E-02     |2.82E-03                   |2.82E-03                  |                             |                            | +/-2.82E-03    | Jy       | 2014ApJS..212...18B |uncertainty                   | 12320   A          | Broad-band measurement                                                                      | 233.73850000 23.50317000 (J2000) |Flux in fixed aperture                                     |  80"x36" aperture                        |From new raw data; Extinction-corrected for Milky Way                                                                                                               
 57     |J (2MASS) AB        |1.2E+01               |+/-0.05      |mag               |2.43E+14  |5.91E-02     |2.72E-03                   |2.72E-03                  |                             |                            | +/-2.72E-03    | Jy       | 2014ApJS..212...18B |uncertainty                   | 12320   A          | Broad-band measurement                                                                      | 233.73850000 23.50317000 (J2000) |Flux in fixed aperture                                     |  80"x36" aperture                        |From new raw data                                                                                                                                                   
 58     |F_J (total)         |1.9E+00               |+/-1.31      |log milliJy       |2.41E+14  |7.94E-02     |2.06E-02                   |2.06E-02                  |                             |                            | +/-2.06E-02    | Jy       | 1995ApJ...453..616S |1 sigma                       | 1.244      microns | Broad-band measurement                                                                      |                                  |Corrected to total flux from single aperture measurement   |                                          |Homogenized from new and previously published data                                                                                                                  
 59     |J_20 (2MASS LGA)    |1.1E+01               |+/-0.019     |mag               |2.40E+14  |5.22E-02     |9.22E-04                   |9.22E-04                  |                             |                            | +/-9.22E-04    | Jy       | 2003AJ....125..525J |1 sigma uncert.               | 1.25      microns  | Broad-band measurement                                                                      | 153457.27 +233010.5 (J2000)      |Flux integrated from map                                   |  45.0 x   45.0 arcsec integration area.  |From new raw data                                                                                                                                                   
 60     |J_Kron (2MASS LGA)  |1.1E+01               |+/-0.019     |mag               |2.40E+14  |5.22E-02     |9.22E-04                   |9.22E-04                  |                             |                            | +/-9.22E-04    | Jy       | 2003AJ....125..525J |1 sigma uncert.               | 1.25      microns  | Broad-band measurement                                                                      | 153457.27 +233010.5 (J2000)      |Flux integrated from map                                   |  45.0 x   45.0 arcsec integration area.  |From new raw data                                                                                                                                                   
 61     |J_tot (2MASS LGA)   |1.1E+01               |+/-0.026     |mag               |2.40E+14  |6.14E-02     |1.49E-03                   |1.49E-03                  |                             |                            | +/-1.49E-03    | Jy       | 2003AJ....125..525J |1 sigma uncert.               | 1.25      microns  | Broad-band measurement                                                                      | 153457.27 +233010.5 (J2000)      |Total flux                                                 |                                          |From new raw data                                                                                                                                                   
 62     |J_14arcsec (2MASS)  |1.2E+01               |+/-0.017     |mag               |2.40E+14  |2.43E-02     |3.83E-04                   |3.83E-04                  |                             |                            | +/-3.83E-04    | Jy       | 20032MASX.C.......: |1 sigma uncert.               | 1.25      microns  | Broad-band measurement                                                                      | 153457.27 +233010.5 (J2000)      |Flux in fixed aperture                                     |  14.0 x 14.0 arcsec aperture             |From new raw data                                                                                                                                                   
 63     |H (ESO/SPM)         |4.5E+01               |+/-3.00      |milliJy           |1.90E+14  |4.51E-02     |3.00E-03                   |3.00E-03                  |                             |                            | +/-3.00E-03    | Jy       | 1995ApJ...453..616S |rms uncertainty               | 1.580      microns | Broad-band measurement                                                                      | 153246.8 +234007 (B1950)         |Flux in fixed aperture                                     |  15" aperture                            |From new raw data                                                                                                                                                   
 64     |F_H (total)         |2.2E+00               |+/-1.57      |log milliJy       |1.84E+14  |1.45E-01     |3.74E-02                   |3.74E-02                  |                             |                            | +/-3.74E-02    | Jy       | 1995ApJ...453..616S |1 sigma                       | 1.634      microns | Broad-band measurement                                                                      |                                  |Corrected to total flux from single aperture measurement   |                                          |Homogenized from new and previously published data                                                                                                                  
 65     |H_20 (2MASS LGA)    |1.0E+01               |+/-0.019     |mag               |1.82E+14  |7.00E-02     |1.24E-03                   |1.24E-03                  |                             |                            | +/-1.24E-03    | Jy       | 2003AJ....125..525J |1 sigma uncert.               | 1.65      microns  | Broad-band measurement                                                                      | 153457.27 +233010.5 (J2000)      |Flux integrated from map                                   |  45.0 x   45.0 arcsec integration area.  |From new raw data                                                                                                                                                   
 66     |H_Kron (2MASS LGA)  |1.0E+01               |+/-0.019     |mag               |1.82E+14  |7.01E-02     |1.24E-03                   |1.24E-03                  |                             |                            | +/-1.24E-03    | Jy       | 2003AJ....125..525J |1 sigma uncert.               | 1.65      microns  | Broad-band measurement                                                                      | 153457.27 +233010.5 (J2000)      |Flux integrated from map                                   |  45.0 x   45.0 arcsec integration area.  |From new raw data                                                                                                                                                   
 67     |H (UH)              |1.1E+01               |+/-0.07      |mag               |1.82E+14  |4.42E-02     |2.85E-03                   |2.85E-03                  |                             |                            | +/-2.85E-03    | Jy       | 2000ApJ...529..170S |uncertainty                   | 1.65   microns     | Broad-band measurement                                                                      | 15 34 57.3 +23 30 11.9 (J2000)   |Flux in fixed aperture                                     |                                          |From new raw data                                                                                                                                                   
 68     |H (UH)              |1.2E+01               |+/-0.1       |mag               |1.82E+14  |2.38E-02     |2.19E-03                   |2.19E-03                  |                             |                            | +/-2.19E-03    | Jy       | 2000ApJ...529..170S |uncertainty                   | 1.65   microns     | Broad-band measurement                                                                      | 15 34 57.3 +23 30 11.9 (J2000)   |Flux in fixed aperture                                     |  Nuclear mag                             |From new raw data                                                                                                                                                   
 69     |H_tot (2MASS LGA)   |1.0E+01               |+/-0.028     |mag               |1.82E+14  |7.72E-02     |2.02E-03                   |2.02E-03                  |                             |                            | +/-2.02E-03    | Jy       | 2003AJ....125..525J |1 sigma uncert.               | 1.65      microns  | Broad-band measurement                                                                      | 153457.27 +233010.5 (J2000)      |Total flux                                                 |                                          |From new raw data                                                                                                                                                   
 70     |H_14arcsec (2MASS)  |1.1E+01               |+/-0.017     |mag               |1.82E+14  |3.69E-02     |5.83E-04                   |5.83E-04                  |                             |                            | +/-5.83E-04    | Jy       | 20032MASX.C.......: |1 sigma uncert.               | 1.65      microns  | Broad-band measurement                                                                      | 153457.27 +233010.5 (J2000)      |Flux in fixed aperture                                     |  14.0 x 14.0 arcsec aperture             |From new raw data                                                                                                                                                   
 71     |H (2MASS) AB        |1.2E+01               |+/-0.06      |mag               |1.82E+14  |7.37E-02     |4.09E-03                   |4.09E-03                  |                             |                            | +/-4.09E-03    | Jy       | 2014ApJS..212...18B |uncertainty                   | 16440   A          | Broad-band measurement                                                                      | 233.73850000 23.50317000 (J2000) |Flux in fixed aperture                                     |  80"x36" aperture                        |From new raw data; Extinction-corrected for Milky Way                                                                                                               
 72     |H (2MASS) AB        |1.2E+01               |+/-0.06      |mag               |1.82E+14  |7.20E-02     |4.00E-03                   |4.00E-03                  |                             |                            | +/-4.00E-03    | Jy       | 2014ApJS..212...18B |uncertainty                   | 16440   A          | Broad-band measurement                                                                      | 233.73850000 23.50317000 (J2000) |Flux in fixed aperture                                     |  80"x36" aperture                        |From new raw data                                                                                                                                                   
 73     |K' (UH)             |1.1E+01               |+/-0.1       |mag               |1.41E+14  |3.10E-02     |2.85E-03                   |2.85E-03                  |                             |                            | +/-2.85E-03    | Jy       | 2000ApJ...529..170S |uncertainty                   | 2.12   microns     | Broad-band measurement                                                                      | 15 34 57.3 +23 30 11.9 (J2000)   |Flux in fixed aperture                                     |  Nuclear mag                             |From new raw data                                                                                                                                                   
 74     |K' (UH)             |1.1E+01               |+/-0.07      |mag               |1.41E+14  |4.01E-02     |2.59E-03                   |2.59E-03                  |                             |                            | +/-2.59E-03    | Jy       | 2000ApJ...529..170S |uncertainty                   | 2.12   microns     | Broad-band measurement                                                                      | 15 34 57.3 +23 30 11.9 (J2000)   |Flux in fixed aperture                                     |                                          |From new raw data                                                                                                                                                   
 75     |Ks (2MASS) AB       |1.2E+01               |+/-0.05      |mag               |1.39E+14  |8.00E-02     |3.68E-03                   |3.68E-03                  |                             |                            | +/-3.68E-03    | Jy       | 2014ApJS..212...18B |uncertainty                   | 21590   A          | Broad-band measurement                                                                      | 233.73850000 23.50317000 (J2000) |Flux in fixed aperture                                     |  80"x36" aperture                        |From new raw data; Extinction-corrected for Milky Way                                                                                                               
 76     |Ks (2MASS) AB       |1.2E+01               |+/-0.05      |mag               |1.39E+14  |7.87E-02     |3.63E-03                   |3.63E-03                  |                             |                            | +/-3.63E-03    | Jy       | 2014ApJS..212...18B |uncertainty                   | 21590   A          | Broad-band measurement                                                                      | 233.73850000 23.50317000 (J2000) |Flux in fixed aperture                                     |  80"x36" aperture                        |From new raw data                                                                                                                                                   
 77     |K_tot (2MASS LGA)   |9.9E+00               |+/-0.036     |mag               |1.38E+14  |7.64E-02     |2.58E-03                   |2.58E-03                  |                             |                            | +/-2.58E-03    | Jy       | 2003AJ....125..525J |1 sigma uncert.               | 2.17      microns  | Broad-band measurement                                                                      | 153457.27 +233010.5 (J2000)      |Total flux                                                 |                                          |From new raw data                                                                                                                                                   
 78     |K_Kron (2MASS LGA)  |1.0E+01               |+/-0.023     |mag               |1.38E+14  |6.94E-02     |1.49E-03                   |1.49E-03                  |                             |                            | +/-1.49E-03    | Jy       | 2003AJ....125..525J |1 sigma uncert.               | 2.17      microns  | Broad-band measurement                                                                      | 153457.27 +233010.5 (J2000)      |Flux integrated from map                                   |  45.0 x   45.0 arcsec integration area.  |From new raw data                                                                                                                                                   
 79     |K_s_14arcsec (2MASS)|1.1E+01               |+/-0.018     |mag               |1.38E+14  |4.03E-02     |6.73E-04                   |6.73E-04                  |                             |                            | +/-6.73E-04    | Jy       | 20032MASX.C.......: |1 sigma uncert.               | 2.17      microns  | Broad-band measurement                                                                      | 153457.27 +233010.5 (J2000)      |Flux in fixed aperture                                     |  14.0 x 14.0 arcsec aperture             |From new raw data                                                                                                                                                   
 80     |K_20 (2MASS LGA)    |1.0E+01               |+/-0.023     |mag               |1.38E+14  |6.94E-02     |1.49E-03                   |1.49E-03                  |                             |                            | +/-1.49E-03    | Jy       | 2003AJ....125..525J |1 sigma uncert.               | 2.17      microns  | Broad-band measurement                                                                      | 153457.27 +233010.5 (J2000)      |Flux integrated from map                                   |  45.0 x   45.0 arcsec integration area.  |From new raw data                                                                                                                                                   
 81     |F_K (total)         |2.1E+00               |+/-1.50      |log milliJy       |1.37E+14  |1.23E-01     |3.19E-02                   |3.19E-02                  |                             |                            | +/-3.19E-02    | Jy       | 1995ApJ...453..616S |1 sigma                       | 2.194      microns | Broad-band measurement                                                                      |                                  |Corrected to total flux from single aperture measurement   |                                          |Homogenized from new and previously published data                                                                                                                  
 82     |K (ESO/SPM)         |4.1E+01               |+/-2.76      |milliJy           |1.36E+14  |4.14E-02     |2.76E-03                   |2.76E-03                  |                             |                            | +/-2.76E-03    | Jy       | 1995ApJ...453..616S |rms uncertainty               | 2.210      microns | Broad-band measurement                                                                      | 153246.8 +234007 (B1950)         |Flux in fixed aperture                                     |  15" aperture                            |From new raw data                                                                                                                                                   
 86     |3.4 microns WISE AB |1.2E+01               |+/-0.10      |mag               |8.93E+13  |4.36E-02     |4.02E-03                   |4.02E-03                  |                             |                            | +/-4.02E-03    | Jy       | 2014ApJS..212...18B |uncertainty                   | 33570   A          | Broad-band measurement                                                                      | 233.73850000 23.50317000 (J2000) |Flux in fixed aperture                                     |  80"x36" aperture; PSF corr              |From new raw data; Extinction-corrected for Milky Way                                                                                                               
 87     |3.4 microns WISE AB |1.2E+01               |+/-0.10      |mag               |8.93E+13  |4.32E-02     |3.98E-03                   |3.98E-03                  |                             |                            | +/-3.98E-03    | Jy       | 2014ApJS..212...18B |uncertainty                   | 33570   A          | Broad-band measurement                                                                      | 233.73850000 23.50317000 (J2000) |Flux in fixed aperture                                     |  80"x36" aperture; PSF corr              |From new raw data                                                                                                                                                   
 88     |3.6 microns IRAC AB |1.2E+01               |+/-0.10      |mag               |8.46E+13  |4.53E-02     |4.17E-03                   |4.17E-03                  |                             |                            | +/-4.17E-03    | Jy       | 2014ApJS..212...18B |uncertainty                   | 35440   A          | Broad-band measurement                                                                      | 233.73850000 23.50317000 (J2000) |Flux in fixed aperture                                     |  80"x36" aperture                        |From new raw data                                                                                                                                                   
 89     |3.6 microns IRAC AB |1.2E+01               |+/-0.10      |mag               |8.46E+13  |4.57E-02     |4.21E-03                   |4.21E-03                  |                             |                            | +/-4.21E-03    | Jy       | 2014ApJS..212...18B |uncertainty                   | 35440   A          | Broad-band measurement                                                                      | 233.73850000 23.50317000 (J2000) |Flux in fixed aperture                                     |  80"x36" aperture                        |From new raw data; Extinction-corrected for Milky Way                                                                                                               
 92     |4.5 microns IRAC AB |1.2E+01               |+/-0.10      |mag               |6.68E+13  |4.15E-02     |3.82E-03                   |3.82E-03                  |                             |                            | +/-3.82E-03    | Jy       | 2014ApJS..212...18B |uncertainty                   | 44870   A          | Broad-band measurement                                                                      | 233.73850000 23.50317000 (J2000) |Flux in fixed aperture                                     |  80"x36" aperture                        |From new raw data                                                                                                                                                   
 93     |4.5 microns IRAC AB |1.2E+01               |+/-0.10      |mag               |6.68E+13  |4.18E-02     |3.85E-03                   |3.85E-03                  |                             |                            | +/-3.85E-03    | Jy       | 2014ApJS..212...18B |uncertainty                   | 44870   A          | Broad-band measurement                                                                      | 233.73850000 23.50317000 (J2000) |Flux in fixed aperture                                     |  80"x36" aperture                        |From new raw data; Extinction-corrected for Milky Way                                                                                                               
 94     |4.6 microns WISE AB |1.2E+01               |+/-0.10      |mag               |6.51E+13  |3.89E-02     |3.58E-03                   |3.58E-03                  |                             |                            | +/-3.58E-03    | Jy       | 2014ApJS..212...18B |uncertainty                   | 46060   A          | Broad-band measurement                                                                      | 233.73850000 23.50317000 (J2000) |Flux in fixed aperture                                     |  80"x36" aperture; PSF corr              |From new raw data                                                                                                                                                   
 95     |4.6 microns WISE AB |1.2E+01               |+/-0.10      |mag               |6.51E+13  |3.91E-02     |3.60E-03                   |3.60E-03                  |                             |                            | +/-3.60E-03    | Jy       | 2014ApJS..212...18B |uncertainty                   | 46060   A          | Broad-band measurement                                                                      | 233.73850000 23.50317000 (J2000) |Flux in fixed aperture                                     |  80"x36" aperture; PSF corr              |From new raw data; Extinction-corrected for Milky Way                                                                                                               
 97     |5.8 microns IRAC AB |1.1E+01               |+/-0.10      |mag               |5.25E+13  |1.13E-01     |1.04E-02                   |1.04E-02                  |                             |                            | +/-1.04E-02    | Jy       | 2014ApJS..212...18B |uncertainty                   | 57100   A          | Broad-band measurement                                                                      | 233.73850000 23.50317000 (J2000) |Flux in fixed aperture                                     |  80"x36" aperture                        |From new raw data                                                                                                                                                   
 98     |5.8 microns IRAC AB |1.1E+01               |+/-0.10      |mag               |5.25E+13  |1.14E-01     |1.05E-02                   |1.05E-02                  |                             |                            | +/-1.05E-02    | Jy       | 2014ApJS..212...18B |uncertainty                   | 57100   A          | Broad-band measurement                                                                      | 233.73850000 23.50317000 (J2000) |Flux in fixed aperture                                     |  80"x36" aperture                        |From new raw data; Extinction-corrected for Milky Way                                                                                                               
 99     |6 microns (Spitzer) |6.9E+01               |             |milliJy           |5.00E+13  |6.93E-02     |                           |                          |                             |                            |                | Jy       | 2009ApJS..182..628V |no uncertainty reported       | 6 microns          | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  From IRS spectra with 3.3% bandpass     |From new raw data                                                                                                                                                   
 103    |LW2 (ISOCAM)        |1.9E+02               |+/-10        |milliJy           |4.44E+13  |1.91E-01     |1.91E-02                   |1.91E-02                  |                             |                            | +/-1.91E-02    | Jy       | 2004A&A...419..501F |estimated error               | 6.75   microns     | Broad-band measurement                                                                      |                                  |Flux in fixed aperture                                     |  2." diameter aperture                   |From reprocessed raw data                                                                                                                                           
 104    |8.0 microns IRAC AB |1.0E+01               |+/-0.10      |mag               |3.82E+13  |3.14E-01     |2.89E-02                   |2.89E-02                  |                             |                            | +/-2.89E-02    | Jy       | 2014ApJS..212...18B |uncertainty                   | 78410   A          | Broad-band measurement                                                                      | 233.73850000 23.50317000 (J2000) |Flux in fixed aperture                                     |  80"x36" aperture                        |From new raw data                                                                                                                                                   
 105    |8.0 microns IRAC AB |1.0E+01               |+/-0.10      |mag               |3.82E+13  |3.15E-01     |2.90E-02                   |2.90E-02                  |                             |                            | +/-2.90E-02    | Jy       | 2014ApJS..212...18B |uncertainty                   | 78410   A          | Broad-band measurement                                                                      | 233.73850000 23.50317000 (J2000) |Flux in fixed aperture                                     |  80"x36" aperture                        |From new raw data; Extinction-corrected for Milky Way                                                                                                               
 106    |7.9 microns Spitzer |5.8E+02               |             |milliJy           |3.79E+13  |5.82E-01     |                           |                          |                             |                            |                | Jy       | 2011ApJ...730...19S |no uncertainty reported       | 7.9 microns        | Broad-band measurement                                                                      | 15 34 57.24 +23 30 11.7 (J2000)  |Flux integrated from map                                   |                                          |From reprocessed raw data                                                                                                                                           
 107    |8 microns (Spitzer) |5.0E+02               |+/-5   %     |milliJy           |3.75E+13  |5.00E-01     |2.50E-02                   |2.50E-02                  |                             |                            | +/-2.50E-02    | Jy       | 2009ApJ...698.1682W |typical accuracy              | 8 microns          | Broad-band measurement                                                                      | 15 34 57.10 +23 30 11.0 (J2000)  |Peak flux                                                  |                                          |From reprocessed raw data                                                                                                                                           
 110    |10 microns (ISO)    |1.5E-01               |+/-30  %     |Jy                |3.00E+13  |1.47E-01     |4.41E-02                   |4.41E-02                  |                             |                            | +/-4.41E-02    | Jy       | 2001A&A...379..823K |uncertainty                   | 10         microns | Broad-band measurement                                                                      |                                  |Flux in fixed aperture                                     |  Aperture 52"                            |From new raw data                                                                                                                                                   
 113    |10.8 microns MIRLIN |1.4E+02               |+/-8         |milliJy           |2.78E+13  |1.42E-01     |8.00E-03                   |8.00E-03                  |                             |                            | +/-8.00E-03    | Jy       | 2004ApJ...605..156G |statistical error             | 10.8   microns     | Broad-band measurement                                                                      |                                  |Flux in fixed aperture                                     |  1.5" diam aperture                      |From new raw data                                                                                                                                                   
 117    |12 microns WISE AB  |9.7E+00               |+/-0.10      |mag               |2.54E+13  |4.96E-01     |4.57E-02                   |4.57E-02                  |                             |                            | +/-4.57E-02    | Jy       | 2014ApJS..212...18B |uncertainty                   | 118100   A         | Broad-band measurement                                                                      | 233.73850000 23.50317000 (J2000) |Flux in fixed aperture                                     |  80"x36" aperture; PSF corr              |From new raw data                                                                                                                                                   
 118    |12 microns WISE AB  |9.7E+00               |+/-0.10      |mag               |2.54E+13  |4.97E-01     |4.58E-02                   |4.58E-02                  |                             |                            | +/-4.58E-02    | Jy       | 2014ApJS..212...18B |uncertainty                   | 118100   A         | Broad-band measurement                                                                      | 233.73850000 23.50317000 (J2000) |Flux in fixed aperture                                     |  80"x36" aperture; PSF corr              |From new raw data; Extinction-corrected for Milky Way                                                                                                               
 119    |12 microns (ISO)    |6.0E-01               |+/-30  %     |Jy                |2.52E+13  |6.00E-01     |1.80E-01                   |1.80E-01                  |                             |                            | +/-1.80E-01    | Jy       | 2001A&A...379..823K |uncertainty                   | 12         microns | Broad-band measurement                                                                      |                                  |Flux in fixed aperture                                     |  Aperture 52"                            |From new raw data                                                                                                                                                   
 120    |12 microns (IRAS)   |6.1E-01               |+/-0.021     |Jy                |2.50E+13  |6.10E-01     |2.10E-02                   |2.10E-02                  |                             |                            | +/-2.10E-02    | Jy       | 2003AJ....126.1607S |1 sigma                       | 12   microns       | Broad-band measurement                                                                      | 15 34 57.1 +23 30 10 (J2000)     |Total flux                                                 |  Size, Method, Flag codes: RI;see paper  |From reprocessed raw data                                                                                                                                           
 121    |12 microns (IRAS)   |6.4E-01               |+/-0.029     |Jy                |2.50E+13  |6.40E-01     |2.90E-02                   |2.90E-02                  |                             |                            | +/-2.90E-02    | Jy       | 1989AJ.....98..766S |rms noise                     | 12         microns | Broad-band measurement                                                                      | 153246.3 +234008 (B1950)         |Integrated from scans                                      |  Marginally resolved with 0.77' beam     |From reprocessed raw data                                                                                                                                           
 122    |12 microns (IRAS)   |4.8E-01               |+/-5   %     |Jy                |2.50E+13  |4.84E-01     |2.42E-02                   |2.42E-02                  |                             |                            | +/-2.42E-02    | Jy       | 1990IRASF.C...0000M |uncertainty                   | 12        microns  | Broad-band measurement                                                                      | 153246.8 +234007 (B1950)         |Flux in fixed aperture                                     |  IRAS quality flag = 3                   |From new raw data                                                                                                                                                   
 129    |14 microns (IRS)    |9.3E-01               |             |Jy                |2.14E+13  |9.30E-01     |                           |                          |                             |                            |                | Jy       | 2007ApJ...659..296L |no uncertainty reported       | 14   microns       | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  S/N = 150                               |From reprocessed raw data                                                                                                                                           
 134    |15 microns (Spitzer)|1.1E+03               |             |milliJy           |2.00E+13  |1.12E+00     |                           |                          |                             |                            |                | Jy       | 2009ApJS..182..628V |no uncertainty reported       | 15 microns         | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  From IRS spectra with 3.3% bandpass     |From new raw data                                                                                                                                                   
 135    |LW3 (ISOCAM)        |7.7E+02               |+/-20        |milliJy           |2.00E+13  |7.65E-01     |1.53E-01                   |1.53E-01                  |                             |                            | +/-1.53E-01    | Jy       | 2004A&A...419..501F |estimated error               | 15.0   microns     | Broad-band measurement                                                                      |                                  |Flux in fixed aperture                                     |  2." diameter aperture                   |From reprocessed raw data                                                                                                                                           
 136    |15 microns (ISO)    |1.1E+00               |+/-30  %     |Jy                |1.98E+13  |1.14E+00     |3.42E-01                   |3.42E-01                  |                             |                            | +/-3.42E-01    | Jy       | 2001A&A...379..823K |uncertainty                   | 15         microns | Broad-band measurement                                                                      |                                  |Flux in fixed aperture                                     |  Aperture 52"                            |From new raw data                                                                                                                                                   
 145    |20 microns (Spitzer)|2.1E+03               |             |milliJy           |1.50E+13  |2.15E+00     |                           |                          |                             |                            |                | Jy       | 2009ApJS..182..628V |no uncertainty reported       | 20 microns         | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  From IRS spectra with 3.3% bandpass     |From new raw data                                                                                                                                                   
 146    |22 microns WISE AB  |7.4E+00               |+/-0.10      |mag               |1.35E+13  |3.86E+00     |3.56E-01                   |3.56E-01                  |                             |                            | +/-3.56E-01    | Jy       | 2014ApJS..212...18B |uncertainty                   | 221400   A         | Broad-band measurement                                                                      | 233.73850000 23.50317000 (J2000) |Flux in fixed aperture                                     |  80"x36" aper; PSF and filter curve corr |From new raw data; Extinction-corrected for Milky Way                                                                                                               
 147    |22 microns WISE AB  |7.1E+00               |+/-0.10      |mag               |1.35E+13  |5.04E+00     |4.65E-01                   |4.65E-01                  |                             |                            | +/-4.65E-01    | Jy       | 2014ApJS..212...18B |uncertainty                   | 221400   A         | Broad-band measurement                                                                      | 233.73850000 23.50317000 (J2000) |Flux in fixed aperture                                     |  80"x36" aperture; PSF corr              |From new raw data                                                                                                                                                   
 148    |22 microns WISE AB  |7.4E+00               |+/-0.10      |mag               |1.35E+13  |3.86E+00     |3.55E-01                   |3.55E-01                  |                             |                            | +/-3.55E-01    | Jy       | 2014ApJS..212...18B |uncertainty                   | 221400   A         | Broad-band measurement                                                                      | 233.73850000 23.50317000 (J2000) |Flux in fixed aperture                                     |  80"x36" aper; PSF and filter curve corr |From new raw data                                                                                                                                                   
 149    |22 microns WISE AB  |7.1E+00               |+/-0.10      |mag               |1.35E+13  |5.05E+00     |4.65E-01                   |4.65E-01                  |                             |                            | +/-4.65E-01    | Jy       | 2014ApJS..212...18B |uncertainty                   | 221400   A         | Broad-band measurement                                                                      | 233.73850000 23.50317000 (J2000) |Flux in fixed aperture                                     |  80"x36" aperture; PSF corr              |From new raw data; Extinction-corrected for Milky Way                                                                                                               
 150    |24 microns MIPS AB  |7.0E+00               |+/-0.10      |mag               |1.28E+13  |5.57E+00     |5.13E-01                   |5.13E-01                  |                             |                            | +/-5.13E-01    | Jy       | 2014ApJS..212...18B |uncertainty                   | 235100   A         | Broad-band measurement                                                                      | 233.73850000 23.50317000 (J2000) |Flux in fixed aperture                                     |  80"x36" aperture; PSF corr              |From new raw data                                                                                                                                                   
 151    |24 microns MIPS AB  |7.0E+00               |+/-0.10      |mag               |1.28E+13  |5.57E+00     |5.13E-01                   |5.13E-01                  |                             |                            | +/-5.13E-01    | Jy       | 2014ApJS..212...18B |uncertainty                   | 235100   A         | Broad-band measurement                                                                      | 233.73850000 23.50317000 (J2000) |Flux in fixed aperture                                     |  80"x36" aperture; PSF corr              |From new raw data; Extinction-corrected for Milky Way                                                                                                               
 152    |25 microns (ISO)    |8.3E+00               |+/-30  %     |Jy                |1.26E+13  |8.28E+00     |2.48E+00                   |2.48E+00                  |                             |                            | +/-2.48E+00    | Jy       | 2001A&A...379..823K |uncertainty                   | 25         microns | Broad-band measurement                                                                      |                                  |Flux in fixed aperture                                     |  Aperture 52"                            |From new raw data                                                                                                                                                   
 155    |25 microns (Spitzer)|9.6E+03               |             |milliJy           |1.20E+13  |9.60E+00     |                           |                          |                             |                            |                | Jy       | 2009ApJS..182..628V |no uncertainty reported       | 25 microns         | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  From IRS spectra with 3.3% bandpass     |From new raw data                                                                                                                                                   
 156    |25 microns (Spitzer)|7.0E+00               |             |Jy                |1.20E+13  |6.97E+00     |                           |                          |                             |                            |                | Jy       | 2011ApJ...730...19S |no uncertainty reported       | 25 microns         | Broad-band measurement                                                                      | 15 34 57.24 +23 30 11.7 (J2000)  |Flux in fixed aperture                                     |                                          |From reprocessed raw data                                                                                                                                           
 157    |25 microns (IRAS)   |8.0E+00               |+/-0.034     |Jy                |1.20E+13  |8.00E+00     |3.40E-02                   |3.40E-02                  |                             |                            | +/-3.40E-02    | Jy       | 2003AJ....126.1607S |1 sigma                       | 25   microns       | Broad-band measurement                                                                      | 15 34 57.1 +23 30 10 (J2000)     |Total flux                                                 |  Size, Method, Flag codes: UT;see paper  |From reprocessed raw data                                                                                                                                           
 158    |25 microns (IRAS)   |7.9E+00               |+/-5   %     |Jy                |1.20E+13  |7.91E+00     |2.42E-02                   |2.42E-02                  |                             |                            | +/-2.42E-02    | Jy       | 1990IRASF.C...0000M |uncertainty                   | 25        microns  | Broad-band measurement                                                                      | 153246.8 +234007 (B1950)         |Flux in fixed aperture                                     |  IRAS quality flag = 3                   |From new raw data                                                                                                                                                   
 159    |25 microns (IRAS)   |7.9E+00               |+/-0.038     |Jy                |1.20E+13  |7.92E+00     |3.80E-02                   |3.80E-02                  |                             |                            | +/-3.80E-02    | Jy       | 1989AJ.....98..766S |rms noise                     | 25         microns | Broad-band measurement                                                                      | 153246.3 +234008 (B1950)         |Integrated from scans                                      |  Unresolved with 0.78' beam              |From reprocessed raw data                                                                                                                                           
 164    |30 microns (Spitzer)|2.3E+04               |             |milliJy           |9.99E+12  |2.29E+01     |                           |                          |                             |                            |                | Jy       | 2009ApJS..182..628V |no uncertainty reported       | 30 microns         | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  From IRS spectra with 3.3% bandpass     |From new raw data                                                                                                                                                   
 168    |52 microns (ISO)    |1.2E+02               |+/-10.8      |Jy                |5.77E+12  |1.21E+02     |1.08E+01                   |1.08E+01                  |                             |                            | +/-1.08E+01    | Jy       | 2008ApJS..178..280B |uncertainty                   | 52 microns         | Broad-band measurement                                                                      | 15 34 57.34 +23 30 11.9 (J2000)  |Flux integrated from map                                   |                                          |From new raw data                                                                                                                                                   
 169    |57 microns (ISO)    |1.3E+02               |+/-11.8      |Jy                |5.26E+12  |1.34E+02     |1.18E+01                   |1.18E+01                  |                             |                            | +/-1.18E+01    | Jy       | 2008ApJS..178..280B |uncertainty                   | 57 microns         | Broad-band measurement                                                                      | 15 34 57.34 +23 30 11.9 (J2000)  |Flux integrated from map                                   |                                          |From new raw data                                                                                                                                                   
 170    |60 microns (IRAS)   |1.0E+02               |+/-0.112     |Jy                |5.00E+12  |1.04E+02     |1.12E-01                   |1.12E-01                  |                             |                            | +/-1.12E-01    | Jy       | 2003AJ....126.1607S |1 sigma                       | 60   microns       | Broad-band measurement                                                                      | 15 34 57.1 +23 30 10 (J2000)     |Total flux                                                 |  Size, Method, Flag codes: UT;see paper  |From reprocessed raw data                                                                                                                                           
 171    |60 microns (IRAS)   |1.0E+02               |+/-4   %     |Jy                |5.00E+12  |1.04E+02     |4.15E+00                   |4.15E+00                  |                             |                            | +/-4.15E+00    | Jy       | 1990IRASF.C...0000M |uncertainty                   | 60        microns  | Broad-band measurement                                                                      | 153246.8 +234007 (B1950)         |Flux in fixed aperture                                     |  IRAS quality flag = 3                   |From new raw data                                                                                                                                                   
 172    |60 microns (IRAS)   |1.0E+02               |+/-0.144     |Jy                |5.00E+12  |1.03E+02     |1.44E-01                   |1.44E-01                  |                             |                            | +/-1.44E-01    | Jy       | 1989AJ.....98..766S |rms noise                     | 60         microns | Broad-band measurement                                                                      | 153246.3 +234008 (B1950)         |Integrated from scans                                      |  Unresolved with 1.44' beam              |From reprocessed raw data                                                                                                                                           
 173    |60 microns (ISO)    |1.1E+02               |+/-30  %     |Jy                |4.93E+12  |1.13E+02     |3.40E+01                   |3.40E+01                  |                             |                            | +/-3.40E+01    | Jy       | 2001A&A...379..823K |uncertainty                   | 60         microns | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Aperture 46" x 46"                      |From new raw data                                                                                                                                                   
 174    |63 microns (ISO)    |1.5E+02               |+/-15.0      |Jy                |4.76E+12  |1.48E+02     |1.50E+01                   |1.50E+01                  |                             |                            | +/-1.50E+01    | Jy       | 2008ApJS..178..280B |uncertainty                   | 63 microns         | Broad-band measurement                                                                      | 15 34 57.34 +23 30 11.9 (J2000)  |Flux integrated from map                                   |                                          |From new raw data                                                                                                                                                   
 175    |88 microns (ISO)    |1.5E+02               |+/-18.7      |Jy                |3.41E+12  |1.51E+02     |1.87E+01                   |1.87E+01                  |                             |                            | +/-1.87E+01    | Jy       | 2008ApJS..178..280B |uncertainty                   | 88 microns         | Broad-band measurement                                                                      | 15 34 57.34 +23 30 11.9 (J2000)  |Flux integrated from map                                   |                                          |From new raw data                                                                                                                                                   
 176    |90 microns (ISO)    |1.1E+02               |+/-30  %     |Jy                |3.15E+12  |1.12E+02     |3.35E+01                   |3.35E+01                  |                             |                            | +/-3.35E+01    | Jy       | 2001A&A...379..823K |uncertainty                   | 90         microns | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Aperture 46" x 46"                      |From new raw data                                                                                                                                                   
 177    |100 microns (IRAS)  |1.2E+02               |+/-0.138     |Jy                |3.00E+12  |1.15E+02     |1.38E-01                   |1.38E-01                  |                             |                            | +/-1.38E-01    | Jy       | 2003AJ....126.1607S |1 sigma                       | 100   microns      | Broad-band measurement                                                                      | 15 34 57.1 +23 30 10 (J2000)     |Total flux                                                 |  Size, Method, Flag codes: UT;see paper  |From reprocessed raw data                                                                                                                                           
 178    |100 microns (IRAS)  |1.1E+02               |+/-3   %     |Jy                |3.00E+12  |1.12E+02     |3.37E+00                   |3.37E+00                  |                             |                            | +/-3.37E+00    | Jy       | 1990IRASF.C...0000M |uncertainty                   | 100       microns  | Broad-band measurement                                                                      | 153246.8 +234007 (B1950)         |Flux in fixed aperture                                     |  IRAS quality flag = 2                   |From new raw data                                                                                                                                                   
 179    |100 microns (IRAS)  |1.1E+02               |+/-0.207     |Jy                |3.00E+12  |1.14E+02     |2.07E-01                   |2.07E-01                  |                             |                            | +/-2.07E-01    | Jy       | 1989AJ.....98..766S |rms noise                     | 100        microns | Broad-band measurement                                                                      | 153246.3 +234008 (B1950)         |Integrated from scans                                      |  Unresolved with 2.94' beam              |From reprocessed raw data                                                                                                                                           
 180    |120 microns (ISO)   |1.1E+02               |+/-30  %     |Jy                |2.52E+12  |1.09E+02     |3.27E+01                   |3.27E+01                  |                             |                            | +/-3.27E+01    | Jy       | 2001A&A...379..823K |uncertainty                   | 120        microns | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Aperture 184" x 184"                    |From new raw data                                                                                                                                                   
 181    |120 microns (ISO)   |1.2E+02               |+/-0.20      |Jy                |2.52E+12  |1.17E+02     |2.00E-01                   |2.00E-01                  |                             |                            | +/-2.00E-01    | Jy       | 2002ApJ...572..105S |1 sigma uncert.               | 119.0      microns | Broad-band measurement                                                                      |                                  |From fitting to map                                        |                                          |From new raw data                                                                                                                                                   
 182    |122 microns (ISO)   |1.2E+02               |+/-9.5       |Jy                |2.46E+12  |1.18E+02     |9.50E+00                   |9.50E+00                  |                             |                            | +/-9.50E+00    | Jy       | 2008ApJS..178..280B |uncertainty                   | 122 microns        | Broad-band measurement                                                                      | 15 34 57.34 +23 30 11.9 (J2000)  |Flux integrated from map                                   |                                          |From new raw data                                                                                                                                                   
 183    |145 microns (ISO)   |1.0E+02               |+/-10.1      |Jy                |2.07E+12  |1.00E+02     |1.01E+01                   |1.01E+01                  |                             |                            | +/-1.01E+01    | Jy       | 2008ApJS..178..280B |uncertainty                   | 145 microns        | Broad-band measurement                                                                      | 15 34 57.34 +23 30 11.9 (J2000)  |Flux integrated from map                                   |                                          |From new raw data                                                                                                                                                   
 184    |158 microns (ISO)   |8.5E+01               |+/-8.5       |Jy                |1.90E+12  |8.45E+01     |8.50E+00                   |8.50E+00                  |                             |                            | +/-8.50E+00    | Jy       | 2008ApJS..178..280B |uncertainty                   | 158 microns        | Broad-band measurement                                                                      | 15 34 57.34 +23 30 11.9 (J2000)  |Flux integrated from map                                   |                                          |From new raw data                                                                                                                                                   
 185    |150 microns (ISO)   |8.8E+01               |+/-30  %     |Jy                |1.86E+12  |8.79E+01     |2.64E+01                   |2.64E+01                  |                             |                            | +/-2.64E+01    | Jy       | 2001A&A...379..823K |uncertainty                   | 150        microns | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Aperture 184" x 184"                    |From new raw data                                                                                                                                                   
 186    |150 microns (ISO)   |7.9E+01               |+/-0.27      |Jy                |1.86E+12  |7.94E+01     |2.70E-01                   |2.70E-01                  |                             |                            | +/-2.70E-01    | Jy       | 2002ApJ...572..105S |1 sigma uncert.               | 161.0      microns | Broad-band measurement                                                                      |                                  |From fitting to map                                        |                                          |From new raw data                                                                                                                                                   
 187    |170 microns (ISO)   |7.7E+01               |+/-6.7       |Jy                |1.76E+12  |7.71E+01     |6.70E+00                   |6.70E+00                  |                             |                            | +/-6.70E+00    | Jy       | 2008ApJS..178..280B |uncertainty                   | 170 microns        | Broad-band measurement                                                                      | 15 34 57.34 +23 30 11.9 (J2000)  |Flux integrated from map                                   |                                          |From new raw data                                                                                                                                                   
 188    |170 microns (ISO)   |7.1E+01               |+/-0.10      |Jy                |1.72E+12  |7.14E+01     |1.00E-01                   |1.00E-01                  |                             |                            | +/-1.00E-01    | Jy       | 2002ApJ...572..105S |1 sigma uncert.               | 174.0      microns | Broad-band measurement                                                                      |                                  |From fitting to map                                        |                                          |From new raw data                                                                                                                                                   
 189    |180 microns (ISO)   |6.4E+01               |+/-30  %     |Jy                |1.62E+12  |6.40E+01     |1.92E+01                   |1.92E+01                  |                             |                            | +/-1.92E+01    | Jy       | 2001A&A...379..823K |uncertainty                   | 180        microns | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Aperture 184" x 184"                    |From new raw data                                                                                                                                                   
 190    |180 microns (ISO)   |4.1E+01               |+/-0.100     |Jy                |1.62E+12  |4.11E+01     |1.00E-01                   |1.00E-01                  |                             |                            | +/-1.00E-01    | Jy       | 2002ApJ...572..105S |1 sigma uncert.               | 185.5      microns | Broad-band measurement                                                                      |                                  |From fitting to map                                        |                                          |From new raw data                                                                                                                                                   
 192    |200 microns (ISO)   |5.5E+01               |+/-30  %     |Jy                |1.47E+12  |5.48E+01     |1.64E+01                   |1.64E+01                  |                             |                            | +/-1.64E+01    | Jy       | 2001A&A...379..823K |uncertainty                   | 200        microns | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Aperture 184" x 184"                    |From new raw data                                                                                                                                                   
 193    |200 microns (ISO)   |3.1E+01               |+/-0.30      |Jy                |1.47E+12  |3.12E+01     |3.00E-01                   |3.00E-01                  |                             |                            | +/-3.00E-01    | Jy       | 2002ApJ...572..105S |1 sigma uncert.               | 204.6      microns | Broad-band measurement                                                                      |                                  |From fitting to map                                        |                                          |From new raw data                                                                                                                                                   
 196    |250 microns (SPIRE) |3.0E+01               |+/-1.5       |Jy                |1.20E+12  |3.01E+01     |1.50E+00                   |1.50E+00                  |                             |                            | +/-1.50E+00    | Jy       | 2011ApJ...743...94R |uncertainty                   | 250 microns        | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |                                          |From new raw data                                                                                                                                                   
 197    |250 microns (BLAST) |2.4E+01               |             |Jy                |1.20E+12  |2.42E+01     |                           |                          |                             |                            |                | Jy       | 2008ApJ...681..415T |no uncertainty reported       | 250 microns        | Broad-band measurement                                                                      | 15 34 57.21 +23 30 09.5 (J2000)  |Modelled datum                                             |                                          |Averaged from previously published data                                                                                                                             
 200    |350 microns (SPIRE) |1.2E+01               |+/-0.6       |Jy                |8.57E+11  |1.17E+01     |6.00E-01                   |6.00E-01                  |                             |                            | +/-6.00E-01    | Jy       | 2011ApJ...743...94R |uncertainty                   | 350 microns        | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |                                          |From new raw data                                                                                                                                                   
 201    |350 microns (BLAST) |9.8E+00               |             |Jy                |8.57E+11  |9.80E+00     |                           |                          |                             |                            |                | Jy       | 2008ApJ...681..415T |no uncertainty reported       | 350 microns        | Broad-band measurement                                                                      | 15 34 57.21 +23 30 09.5 (J2000)  |Modelled datum                                             |                                          |Averaged from previously published data                                                                                                                             
 202    |350 microns         |1.2E+01               |+/-1.0       |Jy                |8.57E+11  |1.17E+01     |1.00E+00                   |1.00E+00                  |                             |                            | +/-1.00E+00    | Jy       | 1996MNRAS.278.1049R |based on count statistics only| 350        microns | Broad-band measurement                                                                      | 153457.22 +233011.40 (J2000)     |Flux in fixed aperture                                     |  8" FWHP                                 |From new raw data                                                                                                                                                   
 203    |350 microns         |1.1E+01               |+/-3.3       |Jy                |8.57E+11  |1.05E+01     |3.30E+00                   |3.30E+00                  |                             |                            | +/-3.30E+00    | Jy       | 1989ApJ...339..859E |uncertainty                   | 350   microns      | Broad-band measurement                                                                      |                                  |Flux in fixed aperture                                     |  104" aperture                           |From new raw data                                                                                                                                                   
 204    |350 microns         |9.7E+00               |+/-0.34      |Jy                |8.57E+11  |9.74E+00     |3.40E-01                   |3.40E-01                  |                             |                            | +/-3.40E-01    | Jy       | 1999CIT...T00R....B |1 sigma                       | 350        microns | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |                                          |From new raw data                                                                                                                                                   
 210    |689 GHz (SMA)       |2.5E+00               |+/-0.8       |Jy                |6.89E+11  |2.50E+00     |8.00E-01                   |8.00E-01                  |                             |                            | +/-8.00E-01    | Jy       | 2009ApJ...693...56M |uncertainty                   | 689.13 GHz         | Broad-band measurement                                                                      | 15 34 57.19 +23 30 11.3 (J2000)  |Total flux                                                 |                                          |From new raw data                                                                                                                                                   
 211    |450 microns         |3.0E+00               |+/-1.1       |Jy                |6.67E+11  |3.00E+00     |1.10E+00                   |1.10E+00                  |                             |                            | +/-1.10E+00    | Jy       | 1989ApJ...339..859E |uncertainty                   | 450   microns      | Broad-band measurement                                                                      |                                  |Flux in fixed aperture                                     |  104" aperture                           |From new raw data                                                                                                                                                   
 212    |450 microns (SCUBA) |6.3E+03               |+/-786       |milliJy           |6.66E+11  |6.29E+00     |7.86E-01                   |7.86E-01                  |                             |                            | +/-7.86E-01    | Jy       | 2001MNRAS.327..697D |uncertainty                   | 450   microns      | Broad-band measurement                                                                      | 15 34 57.2 +23 30 11 (J2000)     |Flux integrated from map                                   |                                          |From new raw data                                                                                                                                                   
 213    |500 microns (SPIRE) |3.9E+00               |+/-0.2       |Jy                |6.00E+11  |3.90E+00     |2.00E-01                   |2.00E-01                  |                             |                            | +/-2.00E-01    | Jy       | 2011ApJ...743...94R |uncertainty                   | 500 microns        | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |                                          |From new raw data                                                                                                                                                   
 214    |500 microns (BLAST) |3.9E+00               |             |Jy                |6.00E+11  |3.90E+00     |                           |                          |                             |                            |                | Jy       | 2008ApJ...681..415T |no uncertainty reported       | 500 microns        | Broad-band measurement                                                                      | 15 34 57.21 +23 30 09.5 (J2000)  |Modelled datum                                             |                                          |Averaged from previously published data                                                                                                                             
 220    |800 microns         |8.3E-01               |+/-0.056     |Jy                |3.75E+11  |8.25E-01     |5.60E-02                   |5.60E-02                  |                             |                            | +/-5.60E-02    | Jy       | 1996MNRAS.278.1049R |based on count statistics only| 800        microns | Broad-band measurement                                                                      | 153457.22 +233011.40 (J2000)     |Flux in fixed aperture                                     |  19" FWHP                                |From new raw data                                                                                                                                                   
 221    |800 microns         |1.1E+00               |+/-0.4       |Jy                |3.75E+11  |1.10E+00     |4.00E-01                   |4.00E-01                  |                             |                            | +/-4.00E-01    | Jy       | 1989ApJ...339..859E |uncertainty                   | 800   microns      | Broad-band measurement                                                                      |                                  |Flux in fixed aperture                                     |  104" aperture                           |From new raw data                                                                                                                                                   
 227    |850 microns (SCUBA) |4.6E+02               |+/-46.9      |milliJy           |3.53E+11  |4.56E-01     |4.69E-02                   |4.69E-02                  |                             |                            | +/-4.69E-02    | Jy       | 2004MNRAS.352..673A |uncertainty                   | 850 microns        | Broad-band measurement                                                                      | 15 34 57.22 +23 30 11.61 (J2000) |Flux integrated from map                                   |                                          |From new raw data                                                                                                                                                   
 228    |850 microns (SCUBA) |8.3E+02               |+/-86        |milliJy           |3.53E+11  |8.32E-01     |8.60E-02                   |8.60E-02                  |                             |                            | +/-8.60E-02    | Jy       | 2000MNRAS.315..115D |uncertainty                   | 850       microns  | Broad-band measurement                                                                      | 153457.2 +233011 (J2000)         |Flux integrated from map                                   |                                          |From new raw data; Corrected for contaminating sources                                                                                                              
 231    |0.87 mm (SMA)       |4.9E-01               |+/-10  %     |Jy                |3.45E+11  |4.90E-01     |4.90E-02                   |4.90E-02                  |                             |                            | +/-4.90E-02    | Jy       | 2009ApJ...700L.104S |1 sigma                       | 0.87   mm          | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  West nucleaus flux                      |From new raw data                                                                                                                                                   
 232    |0.87 mm (SMA)       |1.8E-01               |+/-10  %     |Jy                |3.45E+11  |1.80E-01     |1.80E-02                   |1.80E-02                  |                             |                            | +/-1.80E-02    | Jy       | 2009ApJ...700L.104S |1 sigma                       | 0.87   mm          | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  East nucleaus flux                      |From new raw data                                                                                                                                                   
 234    |277 GHz (SMA)       |1.5E+02               |+/-19        |milliJy           |2.77E+11  |1.52E-01     |1.90E-02                   |1.90E-02                  |                             |                            | +/-1.90E-02    | Jy       | 2009A&A...493..481A |uncertainty                   | 277  GHz           | Broad-band measurement                                                                      | 15 34 57.23 +23 30 11.5 (J2000)  |Flux integrated from map                                   |  West nucleus                            |From new raw data                                                                                                                                                   
 235    |277 GHz (SMA)       |5.8E+01               |+/-16        |milliJy           |2.77E+11  |5.76E-02     |1.60E-02                   |1.60E-02                  |                             |                            | +/-1.60E-02    | Jy       | 2009A&A...493..481A |uncertainty                   | 277  GHz           | Broad-band measurement                                                                      | 15 34 57.31 +23 30 11.4 (J2000)  |Flux integrated from map                                   |  East nucleus                            |From new raw data                                                                                                                                                   
 236    |1.1 mm (SMA)        |2.0E-01               |+/-15  %     |Jy                |2.73E+11  |2.00E-01     |3.00E-02                   |3.00E-02                  |                             |                            | +/-3.00E-02    | Jy       | 2009ApJ...700L.104S |1 sigma                       | 1.1    mm          | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  West nucleaus flux                      |From new raw data                                                                                                                                                   
 237    |1.1 mm (SMA)        |3.3E-01               |+/-0.05      |Jy                |2.73E+11  |3.30E-01     |5.00E-02                   |5.00E-02                  |                             |                            | +/-5.00E-02    | Jy       | 2009ApJ...700L.104S |uncertainty                   | 1.1    mm          | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |                                          |From new raw data                                                                                                                                                   
 238    |1100 microns        |3.5E-01               |+/-0.019     |Jy                |2.73E+11  |3.50E-01     |1.90E-02                   |1.90E-02                  |                             |                            | +/-1.90E-02    | Jy       | 1996MNRAS.278.1049R |based on count statistics only| 1100       microns | Broad-band measurement                                                                      | 153457.22 +233011.40 (J2000)     |Flux in fixed aperture                                     |  19" FWHP                                |From new raw data                                                                                                                                                   
 239    |1100 microns        |                      |<0.6         |Jy                |2.73E+11  |             |                           |                          |  6.0E-01                    |                            | <6.00E-01      | Jy       | 1989ApJ...339..859E |3 sigma                       | 1100   microns     | Broad-band measurement                                                                      |                                  |Flux in fixed aperture                                     |  104" aperture                           |From new raw data                                                                                                                                                   
 240    |1.1 mm (SMA)        |7.0E-02               |+/-15  %     |Jy                |2.73E+11  |7.00E-02     |1.05E-02                   |1.05E-02                  |                             |                            | +/-1.05E-02    | Jy       | 2009ApJ...700L.104S |1 sigma                       | 1.1    mm          | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  East nucleaus flux                      |From new raw data                                                                                                                                                   
 244    |240.904 GHz (SMA)   |2.2E+02               |             |milliJy           |2.41E+11  |2.16E-01     |                           |                          |                             |                            |                | Jy       | 2011A&A...527A..36M |no uncertainty reported       | 240.904 GHz        | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Beam = 2.9" x 2.2"; PA = -55deg         |From new raw data                                                                                                                                                   
 245    |1.25 mm             |2.3E-01               |+/-0.01      |Jy                |2.40E+11  |2.26E-01     |1.00E-02                   |1.00E-02                  |                             |                            | +/-1.00E-02    | Jy       | 1992PASP..104.1086C |uncertainty                   | 1.25   mm          | Broad-band measurement                                                                      |                                  |Flux in fixed aperture                                     |  30" aperture                            |From new raw data                                                                                                                                                   
 246    |238.920 GHz (SMA)   |2.1E+02               |             |milliJy           |2.39E+11  |2.05E-01     |                           |                          |                             |                            |                | Jy       | 2011A&A...527A..36M |no uncertainty reported       | 238.920 GHz        | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Beam = 3.1" x 2.4"; PA = -54deg         |From new raw data                                                                                                                                                   
 247    |236.936 GHz (SMA)   |2.0E+02               |             |milliJy           |2.37E+11  |2.04E-01     |                           |                          |                             |                            |                | Jy       | 2011A&A...527A..36M |no uncertainty reported       | 236.936 GHz        | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Beam = 2.9" x 2.4"; PA = -50deg         |From new raw data                                                                                                                                                   
 248    |234.952 GHz (SMA)   |1.8E+02               |             |milliJy           |2.35E+11  |1.77E-01     |                           |                          |                             |                            |                | Jy       | 2011A&A...527A..36M |no uncertainty reported       | 234.952 GHz        | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Beam = 3.7" x 2.8"; PA = -41deg         |From new raw data                                                                                                                                                   
 249    |232.968 GHz (SMA)   |1.5E+02               |             |milliJy           |2.33E+11  |1.53E-01     |                           |                          |                             |                            |                | Jy       | 2011A&A...527A..36M |no uncertainty reported       | 232.968 GHz        | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Beam = 2.9" x 2.4"; PA = -47deg         |From new raw data                                                                                                                                                   
 250    |230.904 GHz (SMA)   |5.0E+02               |             |milliJy           |2.31E+11  |5.03E-01     |                           |                          |                             |                            |                | Jy       | 2011A&A...527A..36M |no uncertainty reported       | 230.904 GHz        | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Beam = 2.9" x 2.3"; PA = -61deg         |From new raw data                                                                                                                                                   
 252    |1.3 mm              |1.8E+00               |+/-0.5       |Jy                |2.31E+11  |1.80E+00     |5.00E-01                   |5.00E-01                  |                             |                            | +/-5.00E-01    | Jy       | 1986A&A...166L...8C |statistical error             | 1.3        A       | Broad-band measurement                                                                      |                                  |Flux in fixed aperture                                     |  1/2 power beamwidth=90"; abs errors 20% |From new raw data                                                                                                                                                   
 253    |1.3 mm (NRAO)       |3.4E-01               |+/-0.08      |Jy                |2.31E+11  |3.40E-01     |8.00E-02                   |8.00E-02                  |                             |                            | +/-8.00E-02    | Jy       | 1987ApJ...318..645T |uncertainty                   | 1.3 mm             | Broad-band measurement                                                                      | 153247.3 +234006 (B1950)         |Not reported in paper                                      |  Beam size = 33"                         |From new raw data                                                                                                                                                   
 255    |228.920 GHz (SMA)   |1.9E+02               |             |milliJy           |2.29E+11  |1.94E-01     |                           |                          |                             |                            |                | Jy       | 2011A&A...527A..36M |no uncertainty reported       | 228.920 GHz        | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Beam = 3.2" x 2.4"; PA = -62deg         |From new raw data                                                                                                                                                   
 256    |226.936 GHz (SMA)   |2.0E+02               |             |milliJy           |2.27E+11  |2.02E-01     |                           |                          |                             |                            |                | Jy       | 2011A&A...527A..36M |no uncertainty reported       | 226.936 GHz        | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Beam = 2.9" x 2.6"; PA = -54deg         |From new raw data                                                                                                                                                   
 257    |226 GHz (SMA)       |1.7E+02               |+/-33        |milliJy           |2.26E+11  |1.67E-01     |3.30E-02                   |3.30E-02                  |                             |                            | +/-3.30E-02    | Jy       | 2009ApJ...693...56M |uncertainty                   | 226.46 GHz         | Broad-band measurement                                                                      | 15 34 57.19 +23 30 11.3 (J2000)  |Total flux                                                 |                                          |From new raw data                                                                                                                                                   
 258    |224.952 GHz (SMA)   |1.7E+02               |             |milliJy           |2.25E+11  |1.65E-01     |                           |                          |                             |                            |                | Jy       | 2011A&A...527A..36M |no uncertainty reported       | 224.952 GHz        | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Beam = 3.6" x 2.9"; PA = -49deg         |From new raw data                                                                                                                                                   
 259    |222.968 GHz (SMA)   |1.5E+02               |             |milliJy           |2.23E+11  |1.45E-01     |                           |                          |                             |                            |                | Jy       | 2011A&A...527A..36M |no uncertainty reported       | 222.968 GHz        | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Beam = 2.9" x 2.6"; PA = -49deg         |From new raw data                                                                                                                                                   
 260    |1350 microns (SCUBA)|2.7E+02               |+/-32.3      |milliJy           |2.22E+11  |2.71E-01     |3.23E-02                   |3.23E-02                  |                             |                            | +/-3.23E-02    | Jy       | 2004MNRAS.352..673A |uncertainty                   | 1350 microns       | Broad-band measurement                                                                      | 15 34 57.22 +23 30 11.61 (J2000) |Flux integrated from map                                   |                                          |From new raw data                                                                                                                                                   
 261    |220.984 GHz (SMA)   |2.2E+02               |             |milliJy           |2.21E+11  |2.18E-01     |                           |                          |                             |                            |                | Jy       | 2011A&A...527A..36M |no uncertainty reported       | 220.984 GHz        | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Beam = 9.5" x 6.7"; PA = +47deg         |From new raw data                                                                                                                                                   
 265    |219.000 GHz (SMA)   |2.6E+02               |             |milliJy           |2.19E+11  |2.55E-01     |                           |                          |                             |                            |                | Jy       | 2011A&A...527A..36M |no uncertainty reported       | 219.000 GHz        | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Beam = 7.3" x 4.8"; PA = +76deg         |From new raw data                                                                                                                                                   
 266    |217.016 GHz (SMA)   |1.8E+02               |             |milliJy           |2.17E+11  |1.78E-01     |                           |                          |                             |                            |                | Jy       | 2011A&A...527A..36M |no uncertainty reported       | 217.016 GHz        | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Beam = 8.4" x 6.1"; PA = +77deg         |From new raw data                                                                                                                                                   
 267    |216 GHz (SMA)       |1.6E+02               |+/-32        |milliJy           |2.16E+11  |1.60E-01     |3.20E-02                   |3.20E-02                  |                             |                            | +/-3.20E-02    | Jy       | 2009ApJ...693...56M |uncertainty                   | 216.46 GHz         | Broad-band measurement                                                                      | 15 34 57.19 +23 30 11.3 (J2000)  |Total flux                                                 |                                          |From new raw data                                                                                                                                                   
 268    |215.032 GHz (SMA)   |1.6E+02               |             |milliJy           |2.15E+11  |1.56E-01     |                           |                          |                             |                            |                | Jy       | 2011A&A...527A..36M |no uncertainty reported       | 215.032 GHz        | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Beam = 8.5" x 7.0"; PA = +77deg         |From new raw data                                                                                                                                                   
 269    |213.048 GHz (SMA)   |1.5E+02               |             |milliJy           |2.13E+11  |1.45E-01     |                           |                          |                             |                            |                | Jy       | 2011A&A...527A..36M |no uncertainty reported       | 213.048 GHz        | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Beam = 3.8" x 2.8"; PA = +82deg         |From new raw data                                                                                                                                                   
 270    |210.984 GHz (SMA)   |1.8E+02               |             |milliJy           |2.11E+11  |1.77E-01     |                           |                          |                             |                            |                | Jy       | 2011A&A...527A..36M |no uncertainty reported       | 210.984 GHz        | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Beam = 10.0" x 6.9; PA = +47deg         |From new raw data                                                                                                                                                   
 271    |209.000 GHz (SMA)   |1.8E+02               |             |milliJy           |2.09E+11  |1.75E-01     |                           |                          |                             |                            |                | Jy       | 2011A&A...527A..36M |no uncertainty reported       | 209.000 GHz        | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Beam = 7.6" x 5.0"; PA = +76deg         |From new raw data                                                                                                                                                   
 272    |207.016 GHz (SMA)   |1.4E+02               |             |milliJy           |2.07E+11  |1.43E-01     |                           |                          |                             |                            |                | Jy       | 2011A&A...527A..36M |no uncertainty reported       | 207.016 GHz        | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Beam = 8.8" x 6.2"; PA = +76deg         |From new raw data                                                                                                                                                   
 273    |205.032 GHz (SMA)   |1.4E+02               |             |milliJy           |2.05E+11  |1.35E-01     |                           |                          |                             |                            |                | Jy       | 2011A&A...527A..36M |no uncertainty reported       | 205.032 GHz        | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Beam = 8.8" x 7.3"; PA = +76deg         |From new raw data                                                                                                                                                   
 274    |203.048 GHz (SMA)   |1.5E+02               |             |milliJy           |2.03E+11  |1.52E-01     |                           |                          |                             |                            |                | Jy       | 2011A&A...527A..36M |no uncertainty reported       | 203.048 GHz        | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Beam = 3.9" x 3.0"; PA = +82deg         |From new raw data                                                                                                                                                   
 275    |H_2O (3_13-2_20) VLA|1.7E+02               |             |milliJy           |1.83E+11  |1.70E-01     |                           |                          |                             |                            |                | Jy       | 2006ApJ...649..635R |no uncertainty reported       | 183.3101   GHz     | Line measurement; flux integrated over line; lines measured in emission                     |                                  |Flux integrated from map                                   |                                          |From new raw data                                                                                                                                                   
 276    |2000 microns (SCUBA)|8.8E+01               |+/-8.8       |milliJy           |1.50E+11  |8.81E-02     |8.80E-03                   |8.80E-03                  |                             |                            | +/-8.80E-03    | Jy       | 2004MNRAS.352..673A |uncertainty                   | 2000 microns       | Broad-band measurement                                                                      | 15 34 57.22 +23 30 11.61 (J2000) |Flux integrated from map                                   |                                          |From new raw data                                                                                                                                                   
 283    |87.34 GHz (NMA)     |3.0E+01               |             |milliJy           |8.73E+10  |3.00E-02     |                           |                          |                             |                            |                | Jy       | 2007AJ....134.2366I |no uncertainty reported       | 87.34 GHz          | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |                                          |From new raw data                                                                                                                                                   
 284    |32.5 GHz (EVLA)     |6.0E+01               |+/-2.5       |milliJy           |3.25E+10  |5.95E-02     |2.50E-03                   |2.50E-03                  |                             |                            | +/-2.50E-03    | Jy       | 2011ApJ...739L..25L |statistical error             | 32.5 GHz           | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |                                          |From new raw data                                                                                                                                                   
 285    |8085 MHz            |1.7E-01               |+/-0.02      |Jy                |8.08E+09  |1.70E-01     |1.58E-02                   |1.58E-02                  |                             |                            | +/-1.58E-02    | Jy       | 1983AJ.....88...20C |rms uncertainty               | 8085       MHz     | Broad-band measurement                                                                      | 153246.90 +2340 8.2 (B1950)      |Flux integrated from map                                   |                                          |From new raw data                                                                                                                                                   
 286    |7.0 GHz (ATA)       |1.9E-01               |+/-0.02      |Jy                |7.00E+09  |1.90E-01     |2.00E-02                   |2.00E-02                  |                             |                            | +/-2.00E-02    | Jy       | 2010ApJ...710.1462W |uncertainty                   | 7.0 GHz            | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Calibrator is 3C 286                    |From new raw data                                                                                                                                                   
 287    |6.7 GHz (ATA)       |2.3E-01               |+/-0.03      |Jy                |6.70E+09  |2.30E-01     |3.00E-02                   |3.00E-02                  |                             |                            | +/-3.00E-02    | Jy       | 2010ApJ...710.1462W |uncertainty                   | 6.7 GHz            | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Calibrator is 3C 286                    |From new raw data                                                                                                                                                   
 288    |6.3 GHz (ATA)       |2.0E-01               |+/-0.01      |Jy                |6.30E+09  |2.00E-01     |1.00E-02                   |1.00E-02                  |                             |                            | +/-1.00E-02    | Jy       | 2010ApJ...710.1462W |uncertainty                   | 6.3 GHz            | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Calibrator is 3C 286                    |From new raw data                                                                                                                                                   
 289    |6.3 GHz (ATA)       |2.0E-01               |+/-0.03      |Jy                |6.30E+09  |2.00E-01     |3.00E-02                   |3.00E-02                  |                             |                            | +/-3.00E-02    | Jy       | 2010ApJ...710.1462W |uncertainty                   | 6.3 GHz            | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Calibrator is 3C 48                     |From new raw data                                                                                                                                                   
 290    |6.2 GHz (ATA)       |2.9E-01               |+/-0.03      |Jy                |6.20E+09  |2.90E-01     |3.00E-02                   |3.00E-02                  |                             |                            | +/-3.00E-02    | Jy       | 2010ApJ...710.1462W |uncertainty                   | 6.2 GHz            | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Calibrator is 3C 286                    |From new raw data                                                                                                                                                   
 291    |6.0 GHz (ATA)       |2.2E-01               |+/-0.01      |Jy                |6.00E+09  |2.20E-01     |1.00E-02                   |1.00E-02                  |                             |                            | +/-1.00E-02    | Jy       | 2010ApJ...710.1462W |uncertainty                   | 6.0 GHz            | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Calibrator is 3C 286                    |From new raw data                                                                                                                                                   
 292    |5.95 GHz (EVLA)     |1.9E+02               |+/-0.08      |milliJy           |5.95E+09  |1.95E-01     |8.00E-05                   |8.00E-05                  |                             |                            | +/-8.00E-05    | Jy       | 2011ApJ...739L..25L |statistical error             | 5.95 GHz           | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |                                          |From new raw data                                                                                                                                                   
 293    |5.7 GHz (ATA)       |2.2E-01               |+/-0.01      |Jy                |5.70E+09  |2.20E-01     |1.00E-02                   |1.00E-02                  |                             |                            | +/-1.00E-02    | Jy       | 2010ApJ...710.1462W |uncertainty                   | 5.7 GHz            | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Calibrator is 3C 286                    |From new raw data                                                                                                                                                   
 294    |5.7 GHz (ATA)       |2.0E-01               |+/-0.02      |Jy                |5.70E+09  |2.00E-01     |2.00E-02                   |2.00E-02                  |                             |                            | +/-2.00E-02    | Jy       | 2010ApJ...710.1462W |uncertainty                   | 5.7 GHz            | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Calibrator is 3C 48                     |From new raw data                                                                                                                                                   
 295    |5.4 GHz (ATA)       |2.4E-01               |+/-0.01      |Jy                |5.40E+09  |2.40E-01     |1.00E-02                   |1.00E-02                  |                             |                            | +/-1.00E-02    | Jy       | 2010ApJ...710.1462W |uncertainty                   | 5.4 GHz            | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Calibrator is 3C 286                    |From new raw data                                                                                                                                                   
 296    |CH_2_NH (Arecibo)   |3.5E+00               |+/-0.22      |milliJy           |5.29E+09  |3.50E-03     |2.20E-04                   |2.20E-04                  |                             |                            | +/-2.20E-04    | Jy       | 2008AJ....136..389S |uncertainty                   | 5286.813 MHz       | Line measurement; flux integrated over line; lines measured in emission                     |                                  |Peak flux                                                  |                                          |From new raw data                                                                                                                                                   
 297    |5.2 GHz (ATA)       |2.3E-01               |+/-0.01      |Jy                |5.20E+09  |2.30E-01     |1.00E-02                   |1.00E-02                  |                             |                            | +/-1.00E-02    | Jy       | 2010ApJ...710.1462W |uncertainty                   | 5.2 GHz            | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Calibrator is 3C 286                    |From new raw data                                                                                                                                                   
 298    |5.0 GHz (ATA)       |2.4E-01               |+/-0.02      |Jy                |5.00E+09  |2.40E-01     |2.00E-02                   |2.00E-02                  |                             |                            | +/-2.00E-02    | Jy       | 2010ApJ...710.1462W |uncertainty                   | 5.0 GHz            | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Calibrator is 3C 48                     |From new raw data                                                                                                                                                   
 299    |5.0 GHz (ATA)       |2.3E-01               |+/-0.01      |Jy                |5.00E+09  |2.30E-01     |1.00E-02                   |1.00E-02                  |                             |                            | +/-1.00E-02    | Jy       | 2010ApJ...710.1462W |uncertainty                   | 5.0 GHz            | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Calibrator is 3C 286                    |From new raw data                                                                                                                                                   
 300    |5000 MHz (NRAO)     |1.9E-01               |+/-0.029     |Jy                |5.00E+09  |1.92E-01     |2.90E-02                   |2.90E-02                  |                             |                            | +/-2.90E-02    | Jy       | 1976ApJS...32..171S |uncertainty                   | 5000 MHz           | Broad-band measurement                                                                      | 15 32 44.2 +23 40 10 (B1950)     |Flux integrated from map                                   |                                          |From new raw data                                                                                                                                                   
 301    |4.85 GHz            |2.1E+02               |+/-15  %     |milliJy           |4.85E+09  |2.08E-01     |3.12E-02                   |3.12E-02                  |                             |                            | +/-3.12E-02    | Jy       | 1991ApJS...75....1B |uncertainty                   | 4.85       GHz     | Broad-band measurement                                                                      | 153247.1 +233945 (B1950)         |Peak flux                                                  |                                          |From new raw data; Corrected for contaminating sources                                                                                                              
 302    |4.85 GHz            |2.0E+02               |+/-27        |milliJy           |4.85E+09  |2.04E-01     |2.70E-02                   |2.70E-02                  |                             |                            | +/-2.70E-02    | Jy       | 1991ApJS...75.1011G |rms noise                     | 4.85       GHz     | Broad-band measurement                                                                      | 153247.1 +233949 (B1950)         |Modelled datum                                             |                                          |From new raw data; Corrected for contaminating sources                                                                                                              
 303    |4830 MHz (NRAO)     |2.2E+02               |             |milliJy           |4.83E+09  |2.24E-01     |                           |                          |                             |                            |                | Jy       | 1990ApJS...72..621L |no uncertainty reported       | 4830   MHz         | Broad-band measurement                                                                      | 15 34 58.4 +23 30 42 (J2000)     |Flux integrated from map                                   |  S/N = 32                                |From new raw data                                                                                                                                                   
 304    |4.8 GHz (VLA)       |1.8E+02               |             |milliJy           |4.80E+09  |1.83E-01     |                           |                          |                             |                            |                | Jy       | 2010ApJ...720..555P |no uncertainty reported       | 4.8 GHz            | Broad-band measurement                                                                      | 15 34 57.25 +23 30 11.41 (J2000) |Flux integrated from map                                   |                                          |From new raw data                                                                                                                                                   
 305    |4.7 GHz (ATA)       |2.6E-01               |+/-0.02      |Jy                |4.70E+09  |2.60E-01     |2.00E-02                   |2.00E-02                  |                             |                            | +/-2.00E-02    | Jy       | 2010ApJ...710.1462W |uncertainty                   | 4.7 GHz            | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Calibrator is 3C 286                    |From new raw data                                                                                                                                                   
 306    |4.6 GHz (ATA)       |2.4E-01               |+/-0.02      |Jy                |4.60E+09  |2.40E-01     |2.00E-02                   |2.00E-02                  |                             |                            | +/-2.00E-02    | Jy       | 2010ApJ...710.1462W |uncertainty                   | 4.6 GHz            | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Calibrator is 3C 286                    |From new raw data                                                                                                                                                   
 307    |4.5 GHz (ATA)       |2.4E-01               |+/-0.02      |Jy                |4.50E+09  |2.40E-01     |2.00E-02                   |2.00E-02                  |                             |                            | +/-2.00E-02    | Jy       | 2010ApJ...710.1462W |uncertainty                   | 4.5 GHz            | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Calibrator is 3C 286                    |From new raw data                                                                                                                                                   
 308    |4.4 GHz (ATA)       |2.3E-01               |+/-0.02      |Jy                |4.40E+09  |2.30E-01     |2.00E-02                   |2.00E-02                  |                             |                            | +/-2.00E-02    | Jy       | 2010ApJ...710.1462W |uncertainty                   | 4.4 GHz            | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Calibrator is 3C 286                    |From new raw data                                                                                                                                                   
 309    |4.3 GHz (ATA)       |2.5E-01               |+/-0.02      |Jy                |4.30E+09  |2.50E-01     |2.00E-02                   |2.00E-02                  |                             |                            | +/-2.00E-02    | Jy       | 2010ApJ...710.1462W |uncertainty                   | 4.3 GHz            | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Calibrator is 3C 286                    |From new raw data                                                                                                                                                   
 310    |3.6 GHz (ATA)       |2.4E-01               |+/-0.01      |Jy                |3.60E+09  |2.40E-01     |1.00E-02                   |1.00E-02                  |                             |                            | +/-1.00E-02    | Jy       | 2010ApJ...710.1462W |uncertainty                   | 3.6 GHz            | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Calibrator is 3C 286                    |From new raw data                                                                                                                                                   
 311    |3.5 GHz (ATA)       |2.7E-01               |+/-0.01      |Jy                |3.50E+09  |2.70E-01     |1.00E-02                   |1.00E-02                  |                             |                            | +/-1.00E-02    | Jy       | 2010ApJ...710.1462W |uncertainty                   | 3.5 GHz            | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Calibrator is 3C 286                    |From new raw data                                                                                                                                                   
 312    |3.4 GHz (ATA)       |2.8E-01               |+/-0.01      |Jy                |3.40E+09  |2.80E-01     |1.00E-02                   |1.00E-02                  |                             |                            | +/-1.00E-02    | Jy       | 2010ApJ...710.1462W |uncertainty                   | 3.4 GHz            | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Calibrator is 3C 286                    |From new raw data                                                                                                                                                   
 313    |3.3 GHz (ATA)       |2.7E-01               |+/-0.01      |Jy                |3.30E+09  |2.70E-01     |1.00E-02                   |1.00E-02                  |                             |                            | +/-1.00E-02    | Jy       | 2010ApJ...710.1462W |uncertainty                   | 3.3 GHz            | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Calibrator is 3C 286                    |From new raw data                                                                                                                                                   
 314    |3.2 GHz (ATA)       |2.7E-01               |+/-0.01      |Jy                |3.20E+09  |2.70E-01     |1.00E-02                   |1.00E-02                  |                             |                            | +/-1.00E-02    | Jy       | 2010ApJ...710.1462W |uncertainty                   | 3.2 GHz            | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Calibrator is 3C 286                    |From new raw data                                                                                                                                                   
 315    |2.9 GHz (ATA)       |2.7E-01               |+/-0.01      |Jy                |2.90E+09  |2.70E-01     |1.00E-02                   |1.00E-02                  |                             |                            | +/-1.00E-02    | Jy       | 2010ApJ...710.1462W |uncertainty                   | 2.9 GHz            | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Calibrator is 3C 286                    |From new raw data                                                                                                                                                   
 316    |2695 MHz (NRAO)     |2.8E-01               |+/-0.022     |Jy                |2.70E+09  |2.79E-01     |2.20E-02                   |2.20E-02                  |                             |                            | +/-2.20E-02    | Jy       | 1976ApJS...32..171S |uncertainty                   | 2695 MHz           | Broad-band measurement                                                                      | 15 32 44.2 +23 40 10 (B1950)     |Flux integrated from map                                   |                                          |From new raw data                                                                                                                                                   
 317    |2695 MHz            |2.6E-01               |+/-0.01      |Jy                |2.70E+09  |2.60E-01     |1.31E-02                   |1.31E-02                  |                             |                            | +/-1.31E-02    | Jy       | 1983AJ.....88...20C |rms uncertainty               | 2695       MHz     | Broad-band measurement                                                                      | 153246.90 +2340 8.2 (B1950)      |Flux integrated from map                                   |                                          |From new raw data                                                                                                                                                   
 318    |2.6 GHz (ATA)       |2.8E-01               |+/-0.01      |Jy                |2.60E+09  |2.80E-01     |1.00E-02                   |1.00E-02                  |                             |                            | +/-1.00E-02    | Jy       | 2010ApJ...710.1462W |uncertainty                   | 2.6 GHz            | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Calibrator is 3C 286                    |From new raw data                                                                                                                                                   
 319    |2.6 GHz (ATA)       |2.8E-01               |+/-0.02      |Jy                |2.60E+09  |2.80E-01     |2.00E-02                   |2.00E-02                  |                             |                            | +/-2.00E-02    | Jy       | 2010ApJ...710.1462W |uncertainty                   | 2.6 GHz            | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Calibrator is 3C 48                     |From new raw data                                                                                                                                                   
 320    |2.5 GHz (ATA)       |2.7E-01               |+/-0.02      |Jy                |2.50E+09  |2.70E-01     |2.00E-02                   |2.00E-02                  |                             |                            | +/-2.00E-02    | Jy       | 2010ApJ...710.1462W |uncertainty                   | 2.5 GHz            | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Calibrator is 3C 48                     |From new raw data                                                                                                                                                   
 321    |2.5 GHz (ATA)       |2.9E-01               |+/-0.01      |Jy                |2.50E+09  |2.90E-01     |1.00E-02                   |1.00E-02                  |                             |                            | +/-1.00E-02    | Jy       | 2010ApJ...710.1462W |uncertainty                   | 2.5 GHz            | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Calibrator is 3C 286                    |From new raw data                                                                                                                                                   
 322    |2380 MHz            |3.1E+02               |+/-16.       |milliJy           |2.38E+09  |3.12E-01     |1.60E-02                   |1.60E-02                  |                             |                            | +/-1.60E-02    | Jy       | 1978ApJS...36...53D |rms uncertainty               | 2380       MHz     | Broad-band measurement; peak value reported                                                 |                                  |Peak flux                                                  |                                          |From new raw data                                                                                                                                                   
 323    |2.0 GHz (ATA)       |3.0E-01               |+/-0.01      |Jy                |2.00E+09  |3.00E-01     |1.00E-02                   |1.00E-02                  |                             |                            | +/-1.00E-02    | Jy       | 2010ApJ...710.1462W |uncertainty                   | 2.0 GHz            | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Calibrator is 3C 286                    |From new raw data                                                                                                                                                   
 324    |1.9 GHz (ATA)       |3.0E-01               |+/-0.01      |Jy                |1.90E+09  |3.00E-01     |1.00E-02                   |1.00E-02                  |                             |                            | +/-1.00E-02    | Jy       | 2010ApJ...710.1462W |uncertainty                   | 1.9 GHz            | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Calibrator is 3C 286                    |From new raw data                                                                                                                                                   
 325    |1.8 GHz (ATA)       |3.1E-01               |+/-0.01      |Jy                |1.80E+09  |3.10E-01     |1.00E-02                   |1.00E-02                  |                             |                            | +/-1.00E-02    | Jy       | 2010ApJ...710.1462W |uncertainty                   | 1.8 GHz            | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Calibrator is 3C 286                    |From new raw data                                                                                                                                                   
 326    |1.7 GHz (ATA)       |3.0E-01               |+/-0.01      |Jy                |1.70E+09  |3.00E-01     |1.00E-02                   |1.00E-02                  |                             |                            | +/-1.00E-02    | Jy       | 2010ApJ...710.1462W |uncertainty                   | 1.7 GHz            | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Calibrator is 3C 286                    |From new raw data                                                                                                                                                   
 327    |1.6 GHz (ATA)       |3.1E-01               |+/-0.03      |Jy                |1.60E+09  |3.10E-01     |3.00E-02                   |3.00E-02                  |                             |                            | +/-3.00E-02    | Jy       | 2010ApJ...710.1462W |uncertainty                   | 1.6 GHz            | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Calibrator is 3C 286                    |From new raw data                                                                                                                                                   
 328    |1.5 GHz (ATA)       |2.6E-01               |+/-0.02      |Jy                |1.50E+09  |2.60E-01     |2.00E-02                   |2.00E-02                  |                             |                            | +/-2.00E-02    | Jy       | 2010ApJ...710.1462W |uncertainty                   | 1.5 GHz            | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Calibrator is 3C 286                    |From new raw data                                                                                                                                                   
 330    |1.4 GHz (VLA)       |3.0E+02               |             |milliJy           |1.42E+09  |2.99E-01     |                           |                          |                             |                            |                | Jy       | 2006A&A...449..559B |no uncertainty reported       | 1.42   GHz         | Broad-band measurement                                                                      | 15 32 46.92 +23 40 07.8 (J2000)  |Total flux                                                 |                                          |From new raw data                                                                                                                                                   
 332    |1.40 GHz            |3.0E+02               |             |milliJy           |1.40E+09  |3.02E-01     |                           |                          |                             |                            |                | Jy       | 1992ApJS...79..331W |no uncertainty reported       | 1.4        GHz     | Broad-band measurement                                                                      | 153247.1 +233945 (B1950)         |Peak flux                                                  |                                          |From new raw data                                                                                                                                                   
 333    |1.4GHz              |3.3E+02               |+/-9.8       |milliJy           |1.40E+09  |3.27E-01     |9.80E-03                   |9.80E-03                  |                             |                            | +/-9.80E-03    | Jy       | 1998AJ....115.1693C |uncertainty                   | 1.40   GHz         | Broad-band measurement                                                                      | 15 34 57.26 +23 30 11.1 (J2000)  |Flux integrated from map                                   |                                          |From new raw data                                                                                                                                                   
 334    |1400 MHz            |3.0E-01               |+/-0.04      |Jy                |1.40E+09  |3.00E-01     |3.55E-02                   |3.55E-02                  |                             |                            | +/-3.55E-02    | Jy       | 1983AJ.....88...20C |rms uncertainty               | 1400       MHz     | Broad-band measurement                                                                      | 153246.90 +2340 8.2 (B1950)      |Flux integrated from map                                   |                                          |From reprocessed raw data                                                                                                                                           
 335    |1.4 GHz (ATA)       |3.2E-01               |+/-0.01      |Jy                |1.40E+09  |3.20E-01     |1.00E-02                   |1.00E-02                  |                             |                            | +/-1.00E-02    | Jy       | 2010ApJ...710.1462W |uncertainty                   | 1.4 GHz            | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Calibrator is 3C 286                    |From new raw data                                                                                                                                                   
 336    |1.4 GHz (VLA)       |3.3E+02               |             |milliJy           |1.40E+09  |3.26E-01     |                           |                          |                             |                            |                | Jy       | 2002AJ....124..675C |no uncertainty reported       | 1.4   GHz          | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |                                          |Averaged from previously published data                                                                                                                             
 337    |1.2 GHz (ATA)       |3.7E-01               |+/-0.02      |Jy                |1.20E+09  |3.70E-01     |2.00E-02                   |2.00E-02                  |                             |                            | +/-2.00E-02    | Jy       | 2010ApJ...710.1462W |uncertainty                   | 1.2 GHz            | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Calibrator is 3C 48                     |From new raw data                                                                                                                                                   
 338    |1.2 GHz (ATA)       |3.3E-01               |+/-0.01      |Jy                |1.20E+09  |3.30E-01     |1.00E-02                   |1.00E-02                  |                             |                            | +/-1.00E-02    | Jy       | 2010ApJ...710.1462W |uncertainty                   | 1.2 GHz            | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Calibrator is 3C 286                    |From new raw data                                                                                                                                                   
 339    |1.1 GHz (ATA)       |3.6E-01               |+/-0.02      |Jy                |1.10E+09  |3.60E-01     |2.00E-02                   |2.00E-02                  |                             |                            | +/-2.00E-02    | Jy       | 2010ApJ...710.1462W |uncertainty                   | 1.1 GHz            | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Calibrator is 3C 48                     |From new raw data                                                                                                                                                   
 340    |1.1 GHz (ATA)       |3.4E-01               |+/-0.01      |Jy                |1.10E+09  |3.40E-01     |1.00E-02                   |1.00E-02                  |                             |                            | +/-1.00E-02    | Jy       | 2010ApJ...710.1462W |uncertainty                   | 1.1 GHz            | Broad-band measurement                                                                      |                                  |Flux integrated from map                                   |  Calibrator is 3C 286                    |From new raw data                                                                                                                                                   
 341    |365 MHz (Texas)     |4.4E-01               |+/-0.026     |Jy                |3.65E+08  |4.35E-01     |2.60E-02                   |2.60E-02                  |                             |                            | +/-2.60E-02    | Jy       | 1996AJ....111.1945D |internal error                | 365        MHz     | Broad-band measurement; obtained by interpolation over frequency                            | 153246.819 234008.06 (B1950)     |Integrated from scans                                      |  Model:P;MFlag:+;EFlag:+;LFlag:+.        |From new raw data                                                                                                                                                   
 342    |151 MHz             |4.5E-01               |+/-18.1%     |Jy                |1.51E+08  |4.50E-01     |8.13E-02                   |8.13E-02                  |                             |                            | +/-8.13E-02    | Jy       | 1996MNRAS.282..779W |estimated error               | 151        MHz     | Broad-band measurement                                                                      | 153246.9 +233952 (B1950)         |Flux integrated from map; Beam filling or dilution correcte|d                                         |From new raw data; Corrected for contaminating sources                                                                                                              
