
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-06-16T17:05:57PDT



Photometric Data for HS 1700+6416:[SSE2005] MD0094

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|U_n (WHT) AB        | 27.72     |+/-0.33 |mag                 |8.33E+14|  2.96E-08|+/-9.08E-09|Jy|2005ApJ...626..698S|estimated error|    0.36   microns   | Broad-band measurement|17 00 42.020 64 11 24.224 (J2000)| Flux integrated from map|                                        |From new raw data; derived from a flux in a different bandand a color
2|G (WHT) AB          | 25.66     |+/-0.22 |mag                 |6.38E+14|  1.98E-07|+/-3.99E-08|Jy|2005ApJ...626..698S|estimated error|    0.47   microns   | Broad-band measurement|17 00 42.020 64 11 24.224 (J2000)| Flux integrated from map|                                        |From new raw data; derived from a flux in a different bandand a color
3|G (WHT)             | 25.66     ||mag                 |6.38E+14|  1.98E-07||Jy|2006ApJ...647..128E|no uncertainty reported|    0.47   microns   | Broad-band measurement|| Flux in fixed aperture|                                        |Averaged from previously published data
4|H{alpha} (Keck II)  | 2.8E-17   |+/-0.3E-17|erg s^-1^ cm^-2^    |4.57E+14|  2.80E+06|+/-3.00E+05|Jy-Hz|2006ApJ...646..107E|uncertainty|    6563   A         | Line measurement; flux integrated over line; lines measured in emission|17 00 42.02 +64 11 24.22 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
5|R (WHT) AB          | 24.72     |+/-0.16 |mag                 |4.41E+14|  4.70E-07|+/-6.92E-08|Jy|2005ApJ...626..698S|estimated error|    0.68   microns   | Broad-band measurement|17 00 42.020 64 11 24.224 (J2000)| Flux integrated from map|                                        |From new raw data
6|J (Hale/WIRC)       | 22.11     ||mag                 |2.40E+14|  2.23E-06||Jy|2006ApJ...646..107E|no uncertainty reported|    1.25   microns   | Broad-band measurement|17 00 42.02 +64 11 24.22 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data; derived from aflux in a different band and a color
7|K_s (Hale/WIRC)     | 19.65     ||mag                 |1.39E+14|  9.25E-06||Jy|2006ApJ...646..107E|no uncertainty reported|    2.15   microns   | Broad-band measurement|17 00 42.02 +64 11 24.22 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data
8|K_s (P200) AB       | 21.39     |+/-0.22 |mag                 |1.39E+14|  1.01E-05|+/-2.04E-06|Jy|2005ApJ...626..698S|estimated error|    2.15   microns   | Broad-band measurement|17 00 42.020 64 11 24.224 (J2000)| Flux integrated from map|                                        |From new raw data; derived from a flux in a different bandand a color
9|3.6 microns IRAC AB | 20.59     |+/-0.08 |mag                 |8.33E+13|  2.11E-05|+/-1.55E-06|Jy|2005ApJ...626..698S|estimated error|     3.6   microns   | Broad-band measurement|17 00 42.020 64 11 24.224 (J2000)| Flux integrated from map|                                        |From new raw data
10|4.5 microns IRAC AB | 20.43     |+/-0.03 |mag                 |6.66E+13|  2.44E-05|+/-6.75E-07|Jy|2005ApJ...626..698S|estimated error|     4.5   microns   | Broad-band measurement|17 00 42.020 64 11 24.224 (J2000)| Flux integrated from map|                                        |From new raw data
11|5.8 microns IRAC AB | 20.35     |+/-0.22 |mag                 |5.17E+13|  2.63E-05|+/-5.33E-06|Jy|2005ApJ...626..698S|estimated error|     5.8   microns   | Broad-band measurement|17 00 42.020 64 11 24.224 (J2000)| Flux integrated from map|                                        |From new raw data
12|8.0 microns IRAC AB | 20.28     |+/-0.14 |mag                 |3.75E+13|  2.81E-05|+/-3.62E-06|Jy|2005ApJ...626..698S|estimated error|     8.0   microns   | Broad-band measurement|17 00 42.020 64 11 24.224 (J2000)| Flux integrated from map|                                        |From new raw data
13|CO(3-2) (PdBI)      ||<0.3       |Jy km/s             |3.46E+11|  6.91E+05|1.04E+05|Jy-Hz|2010Natur.463..781T|3 sigma|   345.998 GHz       | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|                                        |From new raw data
