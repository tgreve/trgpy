
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-06-14T16:49:52PDT



Photometric Data for PKS 1623+26:[SSP2004] BX0528

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|U (KPNO) AB         | 24.52     |+/-0.18|mag          |8.44E+14|  5.650e-07|+/- 1.019e-07|Jy|2006ApJ...653.1004R|no uncertainty reported|    3550   A         | Broad-band measurement|123653.66 +621724.3 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data; derived from aflux in a different band and a color
2|G (WHT)             | 23.81     |+/-0.14|mag          |7.38E+14|  1.08643e-06|+/- 1.495e-07|Jy|2006ApJ...647..128E|no uncertainty reported|    0.47   microns   | Broad-band measurement|| Flux in fixed aperture|                                        |Averaged from previously published data
4|J (Hale/WIRC)       | 21.54     ||mag                 |2.40E+14|  3.78E-06||Jy|2006ApJ...646..107E|no uncertainty reported|    1.25   microns   | Broad-band measurement|16 25 56.44 +26 50 15.44 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data; derived from aflux in a different band and a color
5|F160W (HST) AB      | 22.33     |+/-0.06 |mag         |1.87E+14|  4.25E-06|+/-2.35E-07|Jy|2011ApJ...731...65F|uncertainty|     1.603 microns   | Broad-band measurement|| Flux in fixed aperture|                                        |From new raw data
6|K_s (Hale/WIRC)     | 19.75     ||mag                 |1.39E+14|  8.44E-06||Jy|2006ApJ...646..107E|no uncertainty reported|    2.15   microns   | Broad-band measurement|16 25 56.44 +26 50 15.44 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data
