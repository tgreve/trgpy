

Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2010-09-03T10:19:38PDT



Photometric Data for SMM J163554.2+661225
No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|F435W (HST/ACS) AB      |  27.04   |+/-0.03|mag                 |6.92E+14|  5.55e-08|+/-1.53e-09|Jy|2011ApJ...734..121S|uncertainty|      4333 A         | Broad-band measurement|189.121506 62.179565 (J2000)| Total flux|                                        |From reprocessed raw data
1|F555W (HST/ACS) AB      |  26.53   |+/-0.02|mag                 |5.63E+14|  8.88e-08|+/-1.63e-09|Jy|2011ApJ...734..121S|uncertainty|      4333 A         | Broad-band measurement|189.121506 62.179565 (J2000)| Total flux|                                        |From reprocessed raw data
1|F625W (HST/ACS) AB      |  26.37   |+/-0.01|mag                 |4.80E+14|  1.03e-07|+/-9.47e-10|Jy|2011ApJ...734..121S|uncertainty|      4333 A         | Broad-band measurement|189.121506 62.179565 (J2000)| Total flux|                                        |From reprocessed raw data
2|F850LP (HST/ACS)    |  26.08  |+/-0.04 | mag                |3.17E+14|1.34e-07|+/-4.95e-09|Jy|2008A&A...477...55H|3 sigma|      9445 A         | Broad-band measurement|14 00 57.530 +02 52 49.34 (J2000)| Flux in fixed aperture|                                        |From new raw data
3|HST F110W (WFC)           | 25.69     |+/-0.05 |mag             |2.67195e+14|1.92e-07 |+/-8.86e-09|Jy |2011ApJ...728L...4H|uncertainty|     3.550 microns   | Broad-band measurement|09 03 11.6 +00 39 06 (J2000)| Flux in fixed aperture|                                        |From new raw data
6|F160W (HST/NICMOS)  | 25.08    |+/-0.01| mag                |1.87E+14| 3.37e-07 |+/-3.11e-09|Jy|2007A&A...470..467C|internal error|       1.6 microns   | Broad-band measurement| | From fitting to map|                                        |From new raw data
21|450 microns (SCUBA) | 46.4      |+/-13.9 |milliJy             |6.66E+11|  46.4E-03|+/-13.9E-03|Jy|2006MNRAS.368..487K|uncertainty|     450   microns   | Broad-band measurement|163554.2 +661225 (J2000)| Flux integrated from map|                                        |From new raw data
25|850 microns (SCUBA) | 15.9      |+/-0.7  |milliJy             |3.53E+11|  15.9E-03|+/-0.7E-03|Jy|2006MNRAS.368..487K|uncertainty|     850   microns   | Broad-band measurement|163554.2 +661225 (J2000)| Flux integrated from map|                                        |From new raw data
25|850 microns (SCUBA) | 17        |+/-2    |milliJy             |3.53E+11|  17.0E-03|+/-2.0E-03|Jy|2006MNRAS.368..487K|uncertainty|     850   microns   | Broad-band measurement|163554.2 +661225 (J2000)| Flux integrated from map|                                        |From new raw data
