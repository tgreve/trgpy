
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-05-28T01:42:09PDT



Photometric Data for SSA22-LAB18, z=3.090

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|3.6 microns (IRAC)  | 7.3       |+/-0.2  | microJy            |8.44E+13|  7.30E-06|+/-2.00E-07|Jy|2009ApJ...692.1561W|uncertainty|     3.550 microns   | Broad-band measurement|22 17 29.0 +00 07 50.2 (J2000)| Corrected to total flux from single aperture measurement|                                        |From new raw data
2|4.5 microns (IRAC)  | 8.7       |+/-0.3  | microJy            |6.67E+13|  8.70E-06|+/-3.00E-07|Jy|2009ApJ...692.1561W|uncertainty|     4.493 microns   | Broad-band measurement|22 17 29.0 +00 07 50.2 (J2000)| Corrected to total flux from single aperture measurement|                                        |From new raw data
3|4.5 microns (IRAC)  | 8.4       |+/-0.3  |microJy             |6.67E+13|  8.40E-06|+/-3.00E-07|Jy|2011ApJ...728...59C|uncertainty|     4.493 microns   | Broad-band measurement|| Flux in fixed aperture|                                        |From reprocessed raw data
4|5.8 microns (IRAC)  | 15.7      |+/-1.5  | microJy            |5.23E+13|  1.57E-05|+/-1.50E-06|Jy|2009ApJ...692.1561W|uncertainty|     5.731 microns   | Broad-band measurement|22 17 29.0 +00 07 50.2 (J2000)| Corrected to total flux from single aperture measurement|                                        |From new raw data
5|8.0 microns (IRAC)  | 19.2      |+/-1.6  | microJy            |3.81E+13|  1.92E-05|+/-1.60E-06|Jy|2009ApJ...692.1561W|uncertainty|     7.872 microns   | Broad-band measurement|22 17 29.0 +00 07 50.2 (J2000)| Corrected to total flux from single aperture measurement|                                        |From new raw data
6|8.0 microns (IRAC)  | 21.2      |+/-2.4  |microJy             |3.81E+13|  2.12E-05|+/-2.40E-06|Jy|2011ApJ...728...59C|uncertainty|     7.872 microns   | Broad-band measurement|| Flux in fixed aperture|                                        |From reprocessed raw data
7|24 microns (MIPS)   | 123.8     |+/-10.6 | microJy            |1.27E+13|  1.24E-04|+/-1.06E-05|Jy|2009ApJ...692.1561W|uncertainty|     23.68 microns   | Broad-band measurement|22 17 29.0 +00 07 50.2 (J2000)| Corrected to total flux from single aperture measurement|                                        |From new raw data
8|24 microns (MIPS)   | 159       |+/-10   |microJy             |1.27E+13|  1.59E-04|+/-1.00E-05|Jy|2011ApJ...728...59C|uncertainty|     23.68 microns   | Broad-band measurement|| Flux integrated from map|                                        |From reprocessed raw data
7|850 microns (SCUBA) | 11.0      |+/-1.5  |milliJy             |3.53E+11|  1.10E-02|+/-1.50E-03|Jy|2005MNRAS.363.1398G|uncertainty|     850   microns   | Broad-band measurement|22 17 28.90 +00 07 51.0 (J2000)| Flux integrated from map|                                        |From new raw data
7|1100 microns (AZTEC) | 2.33      |+/-0.73  |milliJy           |2.73E+11|  2.33E-03|+/-0.73E-03|Jy|2005MNRAS.363.1398G|uncertainty|     850   microns   | Broad-band measurement|22 17 28.90 +00 07 51.0 (J2000)| Flux integrated from map|                                        |From new raw data
1|3500 microns (PdBI)   |        |<0.13   |mJy                 |8.455E10|         |0.13E-03|Jy|2010ApJ...709..210K|3sigma uncertainty|      3500  microns   | Broad-band measurement|16 35 55.67 +66 12 59.51 (J2000)| Flux integrated from map|                                        |From new raw data
