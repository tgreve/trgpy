
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-06-16T17:09:18PDT



Photometric Data for HS 1700+6416:[SSE2005] BX0691

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|U_n (WHT) AB        | 26.21     |+/-0.27 |mag                 |8.33E+14|  1.19E-07|+/-2.94E-08|Jy|2005ApJ...626..698S|estimated error|    0.36   microns   | Broad-band measurement|17 01 05.996 64 12 10.271 (J2000)| Flux integrated from map|                                        |From new raw data; derived from a flux in a different bandand a color
2|G (WHT) AB          | 25.55     |+/-0.19 |mag                 |6.38E+14|  2.19E-07|+/-3.80E-08|Jy|2005ApJ...626..698S|estimated error|    0.47   microns   | Broad-band measurement|17 01 05.996 64 12 10.271 (J2000)| Flux integrated from map|                                        |From new raw data; derived from a flux in a different bandand a color
3|G (WHT)             | 25.55     ||mag                 |6.38E+14|  2.19E-07||Jy|2006ApJ...647..128E|no uncertainty reported|    0.47   microns   | Broad-band measurement|| Flux in fixed aperture|                                        |Averaged from previously published data
4|H{alpha} (Keck II)  | 7.7E-17   |+/-0.3E-17|erg s^-1^ cm^-2^    |4.57E+14|  7.70E+06|+/-3.00E+05|Jy-Hz|2006ApJ...646..107E|uncertainty|    6563   A         | Line measurement; flux integrated over line; lines measured in emission|17 01 06.00 +64 12 10.27 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
5|R (WHT) AB          | 25.33     |+/-0.16 |mag                 |4.41E+14|  2.68E-07|+/-3.95E-08|Jy|2005ApJ...626..698S|estimated error|    0.68   microns   | Broad-band measurement|17 01 05.996 64 12 10.271 (J2000)| Flux integrated from map|                                        |From new raw data
6|J (Hale/WIRC)       | 22.50     ||mag                 |2.40E+14|  1.56E-06||Jy|2006ApJ...646..107E|no uncertainty reported|    1.25   microns   | Broad-band measurement|17 01 06.00 +64 12 10.27 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data; derived from aflux in a different band and a color
7|K_s (Hale/WIRC)     | 20.68     ||mag                 |1.39E+14|  3.58E-06||Jy|2006ApJ...646..107E|no uncertainty reported|    2.15   microns   | Broad-band measurement|17 01 06.00 +64 12 10.27 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data
8|K_s (P200) AB       | 18.87     |+/-0.23 |mag                 |1.39E+14|  1.03E-04|+/-2.21E-05|Jy|2005ApJ...626..698S|estimated error|    2.15   microns   | Broad-band measurement|17 01 05.996 64 12 10.271 (J2000)| Flux integrated from map|                                        |From new raw data; derived from a flux in a different bandand a color
9|3.6 microns IRAC AB | 21.89     |+/-0.10 |mag                 |8.33E+13|  6.37E-06|+/-5.86E-07|Jy|2005ApJ...626..698S|estimated error|     3.6   microns   | Broad-band measurement|17 01 05.996 64 12 10.271 (J2000)| Flux integrated from map|                                        |From new raw data
10|4.5 microns IRAC AB | 21.65     |+/-0.10 |mag                 |6.66E+13|  7.94E-06|+/-7.31E-07|Jy|2005ApJ...626..698S|estimated error|     4.5   microns   | Broad-band measurement|17 01 05.996 64 12 10.271 (J2000)| Flux integrated from map|                                        |From new raw data
11|5.8 microns IRAC AB | 21.44     |+/-0.12 |mag                 |5.17E+13|  9.64E-06|+/-1.06E-06|Jy|2005ApJ...626..698S|estimated error|     5.8   microns   | Broad-band measurement|17 01 05.996 64 12 10.271 (J2000)| Flux integrated from map|                                        |From new raw data
12|8.0 microns IRAC AB | 22.02     |+/-0.27 |mag                 |3.75E+13|  5.65E-06|+/-1.41E-06|Jy|2005ApJ...626..698S|estimated error|     8.0   microns   | Broad-band measurement|17 01 05.996 64 12 10.271 (J2000)| Flux integrated from map|                                        |From new raw data
13|CO(3-2) (PdBI)      ||<0.05      |Jy km/s             |3.46E+11|  5.43E+04|1.81E+04|Jy-Hz|2010Natur.463..781T|3 sigma|   345.998 GHz       | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|                                        |From new raw data
