
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-02-19T10:44:29PST



Photometric Data for AzGN 01

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|U (KPNO) AB         | |>26.7      |mag                 |8.44E+14| |7.59E-08|Jy|2009A&A...500..705M|3 sigma|      3552 A         | Broad-band measurement|12 37 11.9 +62 22 12.4 (J2000)| Flux in fixed aperture|                                        |From new raw data
2|B (HST/ACS) AB          | |>26.3      |mag                 |6.98E+14| |1.10E-07|Jy|2009A&A...500..705M|3 sigma|      4297 A         | Broad-band measurement|12 37 11.9 +62 22 12.4 (J2000)| Flux in fixed aperture|                                        |From new raw data
3|V (HST/ACS) AB          | 25.185    | |mag                 |5.08E+14|  3.06E-07| |Jy|2009A&A...500..705M|no uncertainty reported|      5907 A         | Broad-band measurement|12 37 11.9 +62 22 12.4 (J2000)| Flux in fixed aperture|                                        |From new raw data
4|R (Keck II) AB      | 25.19     | | mag                |4.62E+14|  3.05E-07| |Jy|2004AJ....127.3121W|no uncertainty reported|   648.7   A         | Broad-band measurement|12 37 11.815 +62 22 11.84 (J2000)| Total flux|                                        |From new raw data
5|i (HST/ACS) AB          | 24.487    | |mag                 |3.86E+14|  5.82E-07| |Jy|2009A&A...500..705M|no uncertainty reported|      7764 A         | Broad-band measurement|12 37 11.9 +62 22 12.4 (J2000)| Flux in fixed aperture|                                        |From new raw data
6|z (HST/ACS) AB          | 24.155    | |mag                 |3.17E+14|  7.91E-07| |Jy|2009A&A...500..705M|no uncertainty reported|      9445 A         | Broad-band measurement|12 37 11.9 +62 22 12.4 (J2000)| Flux in fixed aperture|                                        |From new raw data
7|J (KPNO) AB         | |>23.3      |mag                 |2.40E+14| |1.74E-06|Jy|2009A&A...500..705M|3 sigma|  1247.975 nm        | Broad-band measurement|12 37 11.9 +62 22 12.4 (J2000)| Flux in fixed aperture|                                        |From new raw data
8|H (KPNO) AB         | |>23.0      |mag                 |1.83E+14| |2.29E-06|Jy|2009A&A...500..705M|3 sigma|    1635.6 nm        | Broad-band measurement|12 37 11.9 +62 22 12.4 (J2000)| Flux in fixed aperture|                                        |From new raw data
9|K_s(KPNO) AB        | 22.753    | |mag                 |1.40E+14|  2.88E-06| |Jy|2009A&A...500..705M|no uncertainty reported|    2147.5 nm        | Broad-band measurement|12 37 11.9 +62 22 12.4 (J2000)| Flux in fixed aperture|                                        |From new raw data
10|3.6 microns IRAC AB | 21.874    | |mag                 |8.44E+13|  6.46E-06| |Jy|2009A&A...500..705M|no uncertainty reported|     3.550 microns   | Broad-band measurement|12 37 11.9 +62 22 12.4 (J2000)| Flux in fixed aperture|                                        |From new raw data
11|4.5 microns IRAC AB | 21.573    | |mag                 |6.67E+13|  8.53E-06| |Jy|2009A&A...500..705M|no uncertainty reported|     4.493 microns   | Broad-band measurement|12 37 11.9 +62 22 12.4 (J2000)| Flux in fixed aperture|                                        |From new raw data
12|4.5 microns (IRAC)  | 9.5       |+/-1.0  |microJy             |6.67E+13|  9.50E-06|+/-1.00E-06|Jy|2009ApJ...694.1517D|uncertainty|     4.493 microns   | Broad-band measurement|12 37 11.89 +62 22 11.8 (J2000)| Flux integrated from map|                                        |From new raw data
13|5.8 microns IRAC AB | 21.010    | |mag                 |5.23E+13|  1.43E-05| |Jy|2009A&A...500..705M|no uncertainty reported|     5.731 microns   | Broad-band measurement|12 37 11.9 +62 22 12.4 (J2000)| Flux in fixed aperture|                                        |From new raw data
14|8.0 microns IRAC AB | 20.595    | |mag                 |3.81E+13|  2.10E-05| |Jy|2009A&A...500..705M|no uncertainty reported|     7.872 microns   | Broad-band measurement|12 37 11.9 +62 22 12.4 (J2000)| Flux in fixed aperture|                                        |From new raw data
15|8.0 microns (IRAC)  | 26.1      |+/-2.6  |microJy             |3.81E+13|  2.61E-05|+/-2.60E-06|Jy|2009ApJ...694.1517D|uncertainty|     7.872 microns   | Broad-band measurement|12 37 11.89 +62 22 11.8 (J2000)| Flux integrated from map|                                        |From new raw data
17|24 microns (MIPS)   | 65.5      |+/-3.5  |microJy             |1.27E+13|  6.55E-05|+/-3.50E-06|Jy|2009ApJ...694.1517D|uncertainty|     23.68 microns   | Broad-band measurement|12 37 11.89 +62 22 11.8 (J2000)| Flux integrated from map|                                        |From new raw data
18|24 microns (MIPS)   | 68.0      |+/-4.0  |microJy             |1.27E+13|  6.80E-05|+/-4.00E-06|Jy|2009ApJ...694.1517D|uncertainty|     23.68 microns   | Broad-band measurement|12 37 11.89 +62 22 11.8 (J2000)| Flux integrated from map|                                        |From new raw data
19|70 microns (MIPS)   | |<3.0|milliJy             |4.20E+12| |3.0E-3|Jy|2006ApJ...647..L9E|3 sigma|     71.42 microns   | Broad-band measurement| | Flux in fixed aperture|Tentative detection                     |From reprocessed raw data
20|70 microns (PACS)  |           |<2.0    |mJy                 |4.283E+12|         |2.0E-03|Jy|2004MNRAS.354..779G|3sigma uncertainty|      1200 microns   | Broad-band measurement|16 36 55.9 +40 59 12 (J2000)| Flux integrated from map|S/N = 3.66                              |From new raw data
21|100 microns (PACS) | 0.7       |+/-0.4  |mJy             |2.998e+12| 0.7E-03 |+/-0.4E-03 |Jy|2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
22|160 microns (PACS) | 5.4       |+/-1.0  |mJy             |1.874e+12| 5.4E-03 |+/-1.0E-03 |Jy|2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
23|250 microns (SPIRE)| 18.6      |+/-2.7  |mJy                 |1.199e+12| 18.6E-03|+/-2.7e-03 |Jy|2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
24|350 microns (SPIRE)| 41.3      |+/-5.2  |mJy                 |8.565E+11| 41.3E-03|+/-5.2E-03|Jy|2004MNRAS.354..779G|3sigma uncertainty|      1200 microns   | Broad-band measurement|16 36 55.9 +40 59 12 (J2000)| Flux integrated from map|S/N = 3.66                              |From new raw data
25|500 microns (SPIRE)| 39.7      |+/-6.1  |mJy                 |5.996E+11| 39.7E-03|+/-6.1E-03|Jy|2004MNRAS.354..779G|3sigma uncertainty|      1200 microns   | Broad-band measurement|16 36 55.9 +40 59 12 (J2000)| Flux integrated from map|S/N = 3.66                              |From new raw data
26|850 microns (SCUBA) | 20.3      |+/-2.1  |milliJy             |3.53E+11|  2.03E-02|+/-2.10E-03|Jy|2005MNRAS.358..149P|uncertainty|     850   microns   | Broad-band measurement|12 37 11.7 +62 22 12 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
27|1.1mm (AzTEC)       | 11.45     |+/-0.99 |milliJy             |2.73E+11| 11.45E-03|+/-0.99E-03|Jy|2008MNRAS.391..1227P|uncertainty|     850   microns   | Broad-band measurement|12 37 11.7 +62 22 12 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
28|1160 microns (Penner)|10.5      |+/-0.7  |mJy                 |2.58442E+11|10.5E-03|+/-0.7E-03|Jy|2004MNRAS.354..779G|3sigma uncertainty|      1200 microns   | Broad-band measurement|16 36 55.9 +40 59 12 (J2000)| Flux integrated from map|S/N = 3.66                              |From new raw data
29|1.2mm (MAMBO-2)     | 9.3       |+/-0.9  |milliJy             |2.50E+11|  9.3E-03 |+/-0.9E-03 |Jy|2008MNRAS.389..14897P|uncertainty|     850   microns   | Broad-band measurement|12 37 11.7 +62 22 12 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
30|160 GHz (PdBI)      | 1.9       |+/-0.2  | milliJy            |1.60E+11|  1.90E-03|+/-2.00E-04|Jy|2009MNRAS.400..670C|uncertainty|     159.9 GHz       | Broad-band measurement|12 37 11.96 +62 22 12.4 (J2000)| Flux integrated from map|8sigma significance                     |From new raw data
31|137 GHz (PdBI)      | 0.89      |+/-0.15 |milliJy             |1.37E+11|  8.90E-04|+/-1.50E-04|Jy|2010ApJ...714.1407C|uncertainty|       137 GHz       | Broad-band measurement|12 37 11.89 +62 22 11.7 (J2000)| Flux integrated from map|                                        |From new raw data
32|3.3 mm (IRAM)       | 0.33      |+/-0.07 |milliJy             |9.08E+10|  3.30E-04|+/-7.00E-05|Jy|2009ApJ...694.1517D|uncertainty|       3.3 mm        | Broad-band measurement|12 37 11.89 +62 22 11.8 (J2000)| Flux integrated from map|                                        |From new raw data
33|45.6 GHz (VLA)      |           |<65.4|microJy             |4.56E+10| |65.4E-06|Jy|2010ApJ...714.1407C|3 sigma|        43 GHz       | Broad-band measurement|12 37 11.89 +62 22 11.7 (J2000)| Flux integrated from map|                                        |From new raw data
34|45.4 GHz (VLA)      | 0.027     |+/-0.028|mJy             |4.54E+10|0.027E-03|+/-0.028E-03|Jy|2010ApJ...714.1407C|2 sigma|        43 GHz       | Broad-band measurement|12 37 11.89 +62 22 11.7 (J2000)| Flux integrated from map|                                        |From new raw data
35|43 GHz (VLA)        | |<174       |microJy             |4.30E+10| |1.74E-04|Jy|2010ApJ...714.1407C|2 sigma|        43 GHz       | Broad-band measurement|12 37 11.89 +62 22 11.7 (J2000)| Flux integrated from map|                                        |From new raw data
36|23 GHz (VLA)        | |<60        |microJy             |2.30E+10| |6.00E-05|Jy|2010ApJ...714.1407C|2 sigma|        23 GHz       | Broad-band measurement|12 37 11.89 +62 22 11.7 (J2000)| Flux integrated from map|                                        |From new raw data
37|1.4 GHz (VLA)       | 79.3      |+/-13.7 |microJy             |1.40E+09|  7.93E-05|+/-1.37E-05|Jy|2010ApJS..188..178M|uncertainty|       1.4 GHz       | Broad-band measurement|12 37 11.89 +62 22 11.8 (J2000)| Total flux; Beam filling or dilution corrected|Major=2.1"; Minor=0.9"; PA=162 deg      |From new raw data
38|1.4 GHz (VLA)       | 58        |+/-16   | microJy            |1.40E+09|  5.80E-05|+/-1.60E-05|Jy|2006MNRAS.371..963B|1 sigma|       1.4 GHz       | Broad-band measurement|12 37 11.875 +62 22 11.54 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
39|1.4 GHz (VLA)       | 75.8      |+/-7.9  |microJy             |1.40E+09|  7.58E-05|+/-7.90E-06|Jy|2009ApJ...694.1517D|uncertainty|       1.4 GHz       | Broad-band measurement|12 37 11.89 +62 22 11.8 (J2000)| Flux integrated from map|                                        |From new raw data
