
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-07-10T07:28:11PDT



Photometric Data for SBS 1542+541

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|2-10 keV (XMM)      | 1.1E-13   || erg/cm^2^/s        |1.45E+18|  7.59E-09||Jy|2009ApJS..183...17Y|no uncertainty reported|      6.00 keV       | Broad-band measurement|154359.44 +535903.2 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
2|2-10 keV (XMM)      | -13.00    ||log(erg/s/cm^2^)    |1.45E+18|  6.90E-09||Jy|2010A&A...515A...2S|no uncertainty reported|      6.00 keV       | Broad-band measurement|| Modelled datum|                                        |From reprocessed raw data; NED frequency assigned tomid-point of band in keV
3|2-10 keV (XMM)      | -13.0     ||log(erg/s/cm^2^)    |1.45E+18|  6.90E-09||Jy|2008A&A...491..425G|no uncertainty reported|      6.00 keV       | Broad-band measurement|| Modelled datum|                                        |From reprocessed raw data; Extinction-corrected for MilkyWay; NED frequency assigned to mid-point of band in keV
4|0.3-10 keV (XMM)    | -12.889   || log(erg/cm^2^/s)   |1.25E+18|  1.03E-08||Jy|2009ApJ...690.1006F|no uncertainty reported|      5.15 keV       | Broad-band measurement|154359.44 +535903.2 (J2000)| Flux integrated from map|                                        |From reprocessed raw data; NED frequency assigned tomid-point of band in keV
5|0.3-10 keV (XMM)    | 0.2E-12   ||erg cm^-2^ s^-1^    |1.25E+18|  1.60E-08||Jy|2005MNRAS.364..195P|no uncertainty reported|    5.15   keV       | Broad-band measurement|15 43 59.4 +53 59 03.0 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
6|0.5-8 keV (Chandra) | -12.880   || log(erg/cm^2^/s)   |1.03E+18|  1.28E-08||Jy|2009ApJ...690..644G|no uncertainty reported|      4.25 keV       | Broad-band measurement|235.99768 53.984228 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
7|0.5-4.5 keV (XMM)   | -13.05    ||log(erg/cm^2^/s)    |6.05E+17|  1.47E-08||Jy|2011A&A...536A..84V|no uncertainty reported|      2.50 keV       | Broad-band measurement|15 43 59.4 +53 59 02 (J2000)| Flux integrated from map|                                        |Averaged from previously published data; NED frequencyassigned to mid-point of band in keV
8|0.5-2 keV (XMM)     | 5.1E-14   || erg/cm^2^/s        |3.02E+17|  1.69E-08||Jy|2009ApJS..183...17Y|no uncertainty reported|      1.25 keV       | Broad-band measurement|154359.44 +535903.2 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
9|0.5-2 keV (XMM)     | -13.29    ||log(erg/s/cm^2^)    |3.02E+17|  1.70E-08||Jy|2010A&A...515A...2S|no uncertainty reported|      1.25 keV       | Broad-band measurement|| Modelled datum|                                        |From reprocessed raw data; NED frequency assigned tomid-point of band in keV
10|0.5-2 keV (XMM)     | -13.3     ||log(erg/s/cm^2^)    |3.02E+17|  1.66E-08||Jy|2008A&A...491..425G|no uncertainty reported|      1.25 keV       | Broad-band measurement|| Modelled datum|                                        |From reprocessed raw data; Extinction-corrected for MilkyWay; NED frequency assigned to mid-point of band in keV
11|FUV (GALEX) AB      | 20.0996   |+/-0.149518|mag                 |1.95E+15|  3.31E-05|+/-4.56E-06|Jy|2012GASC..C...0000S|uncertainty|1538.6     A         | Broad-band measurement|235.99785361384 53.984065179634 (J2000)| Flux integrated from map|Kron flux in elliptical aperture        |From new raw data
12|FUV (GALEX) AB      | 20.4222   |+/-0.177437|mag                 |1.95E+15|  2.46E-05|+/-4.02E-06|Jy|2012GASC..C...0000S|uncertainty|1538.6     A         | Broad-band measurement|235.99785361384 53.984065179634 (J2000)| Flux in fixed aperture|Flux in 7.5 arcsec diameter aperture    |From new raw data
13|1700 A (SDSS)       | -14.912   ||log(erg/cm^2^/s/A)  |1.76E+15|  1.18E-04||Jy|2011MNRAS.410..860A|no uncertainty reported|      1700 A         | Broad-band measurement|235.997696 +53.984211 (J2000)| Flux integrated from map|                                        |From reprocessed raw data
14|1700 A (SDSS)       | -14.884   ||log(erg/cm^2^/s/A)  |1.76E+15|  1.26E-04||Jy|2011MNRAS.410..860A|no uncertainty reported|      1700 A         | Broad-band measurement|235.997696 +53.984211 (J2000)| Flux integrated from map|                                        |From reprocessed raw data
15|NUV (GALEX) AB      | 19.2063   |+/-0.0551225|mag                 |1.29E+15|  7.54E-05|+/-3.83E-06|Jy|2012GASC..C...0000S|uncertainty|2315.7     A         | Broad-band measurement|235.99785361384 53.984065179634 (J2000)| Flux integrated from map|Kron flux in elliptical aperture        |From new raw data
16|NUV (GALEX) AB      | 19.6095   |+/-0.0692650|mag                 |1.29E+15|  5.20E-05|+/-3.32E-06|Jy|2012GASC..C...0000S|uncertainty|2315.7     A         | Broad-band measurement|235.99785361384 53.984065179634 (J2000)| Flux in fixed aperture|Flux in 7.5 arcsec diameter aperture    |From new raw data
17|u (SDSS Petrosian)AB| 17.652    |+/-0.010|asinh mag           |8.36E+14|  3.28E-04|+/-2.95E-06|Jy|2004SDSS2.C...0000:|based on count statistics only|3585       A         | Broad-band measurement|235.997681 53.984226 (J2000)| Modelled datum|From new raw data
18|u (SDSS PSF) AB     | 17.606    |+/-0.020|asinh mag           |8.36E+14|  3.42E-04|+/-6.29E-06|Jy|2007SDSS6.C...0000:|based on count statistics only|3585       A         | Broad-band measurement|235.9976807164 53.9842276849 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
19|u (SDSS PSF) AB     | 17.606    |+/-0.020|asinh mag           |8.36E+14|  3.42E-04|+/-6.18E-06|Jy|2004SDSS2.C...0000:|based on count statistics only|3585       A         | Broad-band measurement|235.997681 53.984226 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
20|u (SDSS Model) AB   | 17.606    |+/-0.010|asinh mag           |8.36E+14|  3.42E-04|+/-3.12E-06|Jy|2004SDSS2.C...0000:|based on count statistics only|3585       A         | Broad-band measurement|235.997681 53.984226 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
21|u (SDSS CModel) AB  | 17.606    ||asinh mag           |8.36E+14|  3.29E-04||Jy|2004SDSS2.C...0000:|no uncertainty reported|3585       A         | Broad-band measurement|235.997681 53.984226 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
22|g (SDSS PSF) AB     | 16.987    |+/-0.020|asinh mag           |6.17E+14|  5.82E-04|+/-1.07E-05|Jy|2007SDSS6.C...0000:|based on count statistics only|4858       A         | Broad-band measurement|235.9976807164 53.9842276849 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
23|g (SDSS Petrosian)AB| 17.004    |+/-0.003|asinh mag           |6.17E+14|  5.74E-04|+/-1.58E-06|Jy|2004SDSS2.C...0000:|based on count statistics only|4858       A         | Broad-band measurement|235.997681 53.984226 (J2000)| Modelled datum|From new raw data
24|g (SDSS Model) AB   | 16.968    |+/-0.004|asinh mag           |6.17E+14|  5.93E-04|+/-2.44E-06|Jy|2004SDSS2.C...0000:|based on count statistics only|4858       A         | Broad-band measurement|235.997681 53.984226 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
25|g (SDSS PSF) AB     | 16.987    |+/-0.020|asinh mag           |6.17E+14|  5.83E-04|+/-1.09E-05|Jy|2004SDSS2.C...0000:|based on count statistics only|4858       A         | Broad-band measurement|235.997681 53.984226 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
26|g (SDSS CModel) AB  | 16.964    ||asinh mag           |6.17E+14|  5.95E-04||Jy|2004SDSS2.C...0000:|no uncertainty reported|4858       A         | Broad-band measurement|235.997681 53.984226 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
27|V                   | 17.1      |+/-0.1  |mag                 |5.42E+14|  5.26E-04|+/-4.85E-05|Jy|2005MNRAS.358..774B|uncertainty|    5530   A         | Broad-band measurement|| Flux in fixed aperture|                                        |From new raw data; Standard Johnson UBVRI filters assumed
28|r (SDSS PSF) AB     | 17.039    |+/-0.019|asinh mag           |4.77E+14|  5.55E-04|+/-9.72E-06|Jy|2007SDSS6.C...0000:|based on count statistics only|6290       A         | Broad-band measurement|235.9976807164 53.9842276849 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; PETROFAINT - Petrosian radius measured at very low surface brightness; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding; CANONICAL_BAND - this band was primary (usually r);|From new raw data
29|r (SDSS PSF) AB     | 17.039    |+/-0.019|asinh mag           |4.77E+14|  5.55E-04|+/-9.78E-06|Jy|2004SDSS2.C...0000:|based on count statistics only|6290       A         | Broad-band measurement|235.997681 53.984226 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; PETROFAINT - Petrosian radius measured at very low surface brightness; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding; CANONICAL_BAND - this band was primary (usually r);|From new raw data
30|r (SDSS Petrosian)AB| 17.088    |+/-0.004|asinh mag           |4.77E+14|  5.31E-04|+/-1.80E-06|Jy|2004SDSS2.C...0000:|based on count statistics only|6290       A         | Broad-band measurement|235.997681 53.984226 (J2000)| Modelled datum|From new raw data
31|r (SDSS Model) AB   | 17.050    |+/-0.005|asinh mag           |4.77E+14|  5.50E-04|+/-2.51E-06|Jy|2004SDSS2.C...0000:|based on count statistics only|6290       A         | Broad-band measurement|235.997681 53.984226 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; PETROFAINT - Petrosian radius measured at very low surface brightness; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding; CANONICAL_BAND - this band was primary (usually r);|From new raw data
32|r (SDSS CModel) AB  | 17.050    ||asinh mag           |4.77E+14|  5.50E-04||Jy|2004SDSS2.C...0000:|no uncertainty reported|6290       A         | Broad-band measurement|235.997681 53.984226 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; PETROFAINT - Petrosian radius measured at very low surface brightness; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding; CANONICAL_BAND - this band was primary (usually r);|From new raw data
33|R_C                 | 16.9      |+/-0.1  |mag                 |4.68E+14|  5.35E-04|+/-4.93E-05|Jy|2005MNRAS.358..774B|uncertainty|    6400   A         | Broad-band measurement|| Flux in fixed aperture|                                        |From new raw data
34|H{alpha} (TNG)      | 5.2E-14   |+/-20  %|erg/s/cm^2^         |4.57E+14|  5.20E+09|+/-1.04E+09|Jy-Hz|2011A&A...531A.128O|uncertainty|      6563 A         | Line measurement; flux integrated over line; lines measured in emission|15 43 59 +53 59 03 (J2000)| From fitting to map|Broad component flux                    |From new raw data
35|H{alpha} (TNG)      | 2.3E-14   |+/-20  %|erg/s/cm^2^         |4.57E+14|  2.30E+09|+/-4.60E+08|Jy-Hz|2011A&A...531A.128O|uncertainty|      6563 A         | Line measurement; flux integrated over line; lines measured in emission|15 43 59 +53 59 03 (J2000)| From fitting to map|Intermediate component flux             |From new raw data
36|i (SDSS Petrosian)AB| 17.001    |+/-0.004|asinh mag           |3.89E+14|  5.75E-04|+/-2.29E-06|Jy|2004SDSS2.C...0000:|based on count statistics only|7706       A         | Broad-band measurement|235.997681 53.984226 (J2000)| Modelled datum|From new raw data
37|i (SDSS CModel) AB  | 16.958    ||asinh mag           |3.89E+14|  5.98E-04||Jy|2004SDSS2.C...0000:|no uncertainty reported|7706       A         | Broad-band measurement|235.997681 53.984226 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; TOO_LARGE - very large object, poorly determined sky, or bad deblend; ELLIPFAINT - no isophotal fits performed; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
38|i (SDSS PSF) AB     | 16.954    |+/-0.017|asinh mag           |3.89E+14|  6.00E-04|+/-9.40E-06|Jy|2007SDSS6.C...0000:|based on count statistics only|7706       A         | Broad-band measurement|235.9976807164 53.9842276849 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; TOO_LARGE - very large object, poorly determined sky, or bad deblend; ELLIPFAINT - no isophotal fits performed; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
39|i (SDSS PSF) AB     | 16.954    |+/-0.017|asinh mag           |3.89E+14|  6.01E-04|+/-9.31E-06|Jy|2004SDSS2.C...0000:|based on count statistics only|7706       A         | Broad-band measurement|235.997681 53.984226 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; TOO_LARGE - very large object, poorly determined sky, or bad deblend; ELLIPFAINT - no isophotal fits performed; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
40|i (SDSS Model) AB   | 16.958    |+/-0.005|asinh mag           |3.89E+14|  5.98E-04|+/-2.99E-06|Jy|2004SDSS2.C...0000:|based on count statistics only|7706       A         | Broad-band measurement|235.997681 53.984226 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; TOO_LARGE - very large object, poorly determined sky, or bad deblend; ELLIPFAINT - no isophotal fits performed; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
41|z (SDSS PSF) AB     | 16.712    |+/-0.020|asinh mag           |3.25E+14|  7.36E-04|+/-1.38E-05|Jy|2004SDSS2.C...0000:|based on count statistics only|9222       A         | Broad-band measurement|235.997681 53.984226 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; ELLIPFAINT - no isophotal fits performed; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
42|z (SDSS Model) AB   | 16.707    |+/-0.010|asinh mag           |3.25E+14|  7.40E-04|+/-6.75E-06|Jy|2004SDSS2.C...0000:|based on count statistics only|9222       A         | Broad-band measurement|235.997681 53.984226 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; ELLIPFAINT - no isophotal fits performed; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
43|z (SDSS CModel) AB  | 16.701    ||asinh mag           |3.25E+14|  7.58E-04||Jy|2004SDSS2.C...0000:|no uncertainty reported|9222       A         | Broad-band measurement|235.997681 53.984226 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; ELLIPFAINT - no isophotal fits performed; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
44|z (SDSS Petrosian)AB| 16.741    |+/-0.013|asinh mag           |3.25E+14|  7.17E-04|+/-8.38E-06|Jy|2004SDSS2.C...0000:|based on count statistics only|9222       A         | Broad-band measurement|235.997681 53.984226 (J2000)| Modelled datum|From new raw data
45|z (SDSS PSF) AB     | 16.712    |+/-0.020|asinh mag           |3.25E+14|  7.37E-04|+/-1.36E-05|Jy|2007SDSS6.C...0000:|based on count statistics only|9222       A         | Broad-band measurement|235.9976807164 53.9842276849 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; ELLIPFAINT - no isophotal fits performed; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
46|J (2MASS)           | 7.28e-04  || Jy                 |2.40E+14|  7.28E-04||Jy|2008MNRAS.383.1513L|no uncertainty reported|      1.25 microns   | Broad-band measurement|15 43 59.44 +53 59 03.2 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data; Extinction-correctedfor Milky Way
47|H (2MASS)           | 9.21e-04  || Jy                 |1.82E+14|  9.21E-04||Jy|2008MNRAS.383.1513L|no uncertainty reported|      1.65 microns   | Broad-band measurement|15 43 59.44 +53 59 03.2 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data; Extinction-correctedfor Milky Way
48|K_s (2MASS)         | 1.22e-03  || Jy                 |1.38E+14|  1.22E-03||Jy|2008MNRAS.383.1513L|no uncertainty reported|      2.17 microns   | Broad-band measurement|15 43 59.44 +53 59 03.2 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data; Extinction-correctedfor Milky Way
49|250 GHz (IRAM/MAMBO)| 3.8E-03   |+/-0.9E-03|Jy                  |2.50E+11|  3.80E-03|+/-9.00E-04|Jy|2006AJ....132.1307P|1 sigma|     250   GHz       | Broad-band measurement|15 43 59.37 +53 59 03.1 (J2000)| Flux integrated from map|From 2003A&A...398..857O                |Averaged from previously published data
49|115GHz              | 0.11E-03   |+/-0.02E-03|Jy                |1.15E+11|  0.11E-03|+/-0.02E-03|Jy|2006AJ....132.1307P|1 sigma|     250   GHz       | Broad-band measurement|15 43 59.37 +53 59 03.1 (J2000)| Flux integrated from map|From 2003A&A...398..857O                |Averaged from previously published data
50|5.0 GHz (VLA)       | 370E-06   |+/-100E-06|Jy                  |5.00E+09|  3.70E-04|+/-1.00E-04|Jy|2006AJ....132.1307P|1 sigma|     5.0   GHz       | Broad-band measurement|15 43 59.37 +53 59 03.1 (J2000)| Flux integrated from map|                                        |From new raw data
51|1.4 GHz (VLA)       | 140E-06   |+/-20E-06|Jy                  |1.40E+09|  1.40E-04|+/-2.00E-05|Jy|2006AJ....132.1307P|1 sigma|     1.4   GHz       | Broad-band measurement|15 43 59.37 +53 59 03.1 (J2000)| Flux integrated from map|                                        |From new raw data
