
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-05-30T01:49:31PDT



Photometric Data for BzK 21000

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
2|3.6 microns (IRAC)  | 40.00     |+/-2.00 |microJy        |8.44E+13|  4.00E-05|+/-2.00E-06|Jy|2011AJ....141....1T|rms uncertainty|     3.550 microns   | Broad-band measurement|189.294266 62.376274 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
3|4.5 microns (IRAC)  | 47.50     |+/-2.38 |microJy        |6.67E+13|  4.75E-05|+/-2.38E-06|Jy|2011AJ....141....1T|rms uncertainty|     4.493 microns   | Broad-band measurement|189.294266 62.376274 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
4|5.8 microns (IRAC)  | 39.60     |+/-2.11 |microJy        |5.23E+13|  3.96E-05|+/-2.11E-06|Jy|2011AJ....141....1T|rms uncertainty|     5.731 microns   | Broad-band measurement|189.294266 62.376274 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
5|8.0 microns (IRAC)  | 44.20     |+/-2.30 |microJy        |3.81E+13|  4.42E-05|+/-2.30E-06|Jy|2011AJ....141....1T|rms uncertainty|     7.872 microns   | Broad-band measurement|189.294266 62.376274 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
6|16 microns (IRS)    | 240.4     |+/-11.5 |microJy        |1.90E+13|  2.40E-04|+/-1.15E-05|Jy|2011AJ....141....1T|rms uncertainty|      15.8 microns   | Broad-band measurement|189.294266 62.376274 (J2000)| From fitting to map|                                        |From new raw data
7|24 microns (MIPS)   | 386.0     |+/-4.9  |microJy        |1.27E+13|  3.86E-04|+/-4.90E-06|Jy|2011AJ....141....1T|rms uncertainty|     23.68 microns   | Broad-band measurement|189.294266 62.376274 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
8|24 microns (MIPS)   | 383.0     |+/-7.0  |microJy        |1.27E+13|  3.83E-04|+/-7.00E-06|Jy|2011AJ....141....1T|rms uncertainty|     23.68 microns   | Broad-band measurement|189.294266 62.376274 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
9|24 microns (MIPS)   | 382.0     |+/-6.0  |microJy        |1.27E+13|  3.82E-04|+/-6.00E-06|Jy|2011AJ....141....1T|rms uncertainty|     23.68 microns   | Broad-band measurement|189.294266 62.376274 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
10|24 microns (Spitzer)| 227      |+/-39   |microJy        |1.27E+13|  2.27E-04|+/-3.90E-05|Jy|2011ApJ...726...93R|uncertainty|     23.68 microns   | Broad-band measurement|12 37 10.60 +62 22 34.6 (J2000)| Not reported in paper|                                        |Averaged from previously published data
11|70 microns (Spitzer)| 3.9      |+/-0.5  |mJy            |4.20E+12|  3.90E-03|+/-5.00E-04|Jy|2009MNRAS.399..121C|uncertainty|     71.42 microns   | Broad-band measurement|123710.60 +622234.6 (J2000)| Flux integrated from map|                                        |From reprocessed raw data
12|70 microns (Spitzer)| 4.9      |+/-0.7  |mJy            |4.20E+12|  4.90E-03|+/-7.00E-04|Jy|2009MNRAS.399..121C|uncertainty|     71.42 microns   | Broad-band measurement|123710.60 +622234.6 (J2000)| Flux integrated from map|                                        |From reprocessed raw data
13|70 microns (PACS)   | 4.9      |+/-0.7  |mJy            |4.283e+12|  4.9E-03 |+/-0.7E-03 |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
14|100 microns (PACS)  | 8.1      |+/-0.6  |mJy            |2.998e+12|  8.1E-03 |+/-0.6E-03 |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
15|160 microns (PACS)  | 15.1     |+/-1.4  |mJy            |1.874e+12|  15.1E-03|+/-1.4E-03 |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
16|250 microns (SPIRE) | 24.4     |+/-2.5  |mJy            |1.199e+12|  24.4E-03 |+/-2.5e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
17|350 microns (SPIRE) | 20.1     |+/-4.7  |mJy            |8.565e+11|  20.1E-03 |+/-4.7e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
18|500 microns (SPIRE) | 11.6     |+/-7.4  |mJy            |5.996e+11|  11.6E-03 |+/-7.4e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
19|850 microns (SCUBA) |          |<1.8    |mJy            |3.53E+11| |1.80E-03|Jy|2009MNRAS.399..121C|2 sigma|       850 microns   | Broad-band measurement|123710.60 +622234.6 (J2000)| Flux integrated from map|                                        |From new raw data
20|1160 microns (Penner)|         |<2.2    |mJy            |2.58442E+11|       |2.2E-03|Jy|2004MNRAS.354..779G|3sigma uncertainty|      1200 microns   | Broad-band measurement|16 36 55.9 +40 59 12 (J2000)| Flux integrated from map|S/N = 3.66                              |From new raw data
21|1200 microns (MAMBO)|          |<1.8    |mJy            |2.50E+11|  |1.8E-03|Jy|2004MNRAS.354..779G|3sigma uncertainty|      1200 microns   | Broad-band measurement|16 36 55.9 +40 59 12 (J2000)| Flux integrated from map|S/N = 3.66                              |From new raw data
25|43.34 GHz (VLA)     |          |<144.0  |uJy            |43.34E+09|  |144.E-06|Jy|2009MNRAS.399..121C|2rms uncertainty|       1.4 GHz       | Broad-band measurement|123710.60 +622234.6 (J2000)| Flux integrated from map|                                        |From new raw data
26|1.4 GHz (MERLIN)    | 38.3     |+/-10.1 |uJy            |1.40E+09|  3.83E-05|+/-1.01E-05|Jy|2009MNRAS.399..121C|uncertainty|       1.4 GHz       | Broad-band measurement|123710.60 +622234.6 (J2000)| Flux integrated from map|                                        |From new raw data
27|1.4 GHz (VLA)       | 42.8     |+/-6.7  |uJy            |1.40E+09|  4.28E-05|+/-6.70E-06|Jy|2010ApJS..188..178M|uncertainty|       1.4 GHz       | Broad-band measurement|12 37 10.60 +62 22 34.6 (J2000)| Total flux; Beam filling or dilution corrected|Major=0.0"; Minor=0.0"; PA=0 deg        |From new raw data
