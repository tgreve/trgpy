
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-07-10T07:09:01PDT



Photometric Data for B1938+666

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
40|850 microns (SCUBA) | 34.6       |+/-2.0  |milliJy             |3.53E+11|  34.6E-03|+/-2.0E-03|Jy|2005MNRAS.358..149P|uncertainty|     850   microns   | Broad-band measurement|12 36 18.7 +62 15 53 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
15|450 microns (SCUBA) | 126       |+/-22   |milliJy             |6.66E+11|  126.0E-03|+/-22.0E-03|Jy|2010A&A...518L..35I|uncertainty|       450 microns   | Broad-band measurement| | Flux integrated from map|                                        |From new raw data
15|1350 microns (SCUBA) | 14.7       |+/-2   |milliJy             |2.22E+11|  14.7E-03|+/-2.0E-03|Jy|2010A&A...518L..35I|uncertainty|       450 microns   | Broad-band measurement| | Flux integrated from map|                                        |From new raw data
15|114 GHz              | 56.27       |+/-5.63   |milliJy             |1.14E+11|  56.27E-03|+/-5.63E-03|Jy|2010A&A...518L..35I|uncertainty|       450 microns   | Broad-band measurement| | Flux integrated from map|                                        |From new raw data
15|113.0425 GHz         | 17.76       |+/-0.26   |milliJy             |113.0425E+09|  17.76E-03|+/-0.26E-03|Jy|2010A&A...518L..35I|uncertainty|       450 microns   | Broad-band measurement| | Flux integrated from map|                                        |From new raw data
15|75.3638 GHz          | 23.89       |+/-0.32   |milliJy             |75.3638E+09|  23.89E-03|+/-0.32E-03|Jy|2010A&A...518L..35I|uncertainty|       450 microns   | Broad-band measurement| | Flux integrated from map|                                        |From new raw data
