

Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.


queryDateTime:2009-11-03T15:07:35PST






Photometric Data for MIPS8196 (z=2.586)

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
4|R (KPNO)            | 3.108     ||microJy             |4.66E+14|  3.11E-06||Jy|2007ApJ...658..778Y|no uncertainty reported|    6440   A         | Broad-band measurement|171510.28 +600955.2 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data
5|R (Cousins) m_aper  | 22.61     |+/-0.03 |mag                 |4.65E+14|  2.77E-06|+/-7.64E-08|Jy|2004AJ....128....1F|based on count statistics only|6440       A         | Broad-band measurement|171510.200 +600954.97 (J2000)| Flux in fixed aperture|3-arcsecond aperture                    |From new raw data
6|R (Cousins) m_tot   | 22.44     |+/-0.04 |mag                 |4.65E+14|  3.23E-06|+/-1.19E-07|Jy|2004AJ....128....1F|based on count statistics only|6440       A         | Broad-band measurement|171510.200 +600954.97 (J2000)| Total flux|                                        |From new raw data
7|F160W (HST NICMOS)  | 18.68     || mag                |1.86E+14|  3.52E-05||Jy|2008ApJ...680..232D|no uncertainty reported|      1.61 microns   | Broad-band measurement|17 15 10.17 +60 09 54.54 (J2000)| Flux integrated from map|                                        |From new raw data
8|3.6 microns (IRAC)  | 81        |+/-6    | microJy            |8.44E+13|  8.10E-05|+/-6.00E-06|Jy|2007ApJ...664..713S|uncertainty|   3.550   microns   | Broad-band measurement|| Flux in fixed aperture|7.3" diameter aperture                  |From reprocessed raw data
9|3.6 microns (IRAC)  | 106.03    |+/-11.72|microJy             |8.42E+13|  1.06E-04|+/-1.17E-05|Jy|2005ApJS..161...41L|uncertainty|3.56       microns   | Broad-band measurement|171510.18 +600954.5 (J2000)| Flux in fixed aperture|Aperture =       7.59 arcsec.           |From new raw data
10|4.5 microns (IRAC)  | 61        |+/-6    | microJy            |6.67E+13|  6.10E-05|+/-6.00E-06|Jy|2007ApJ...664..713S|uncertainty|   4.493   microns   | Broad-band measurement|| Flux in fixed aperture|7.3" diameter aperture                  |From reprocessed raw data
11|4.5 microns (IRAC)  | 89.19     |+/-10.38|microJy             |6.63E+13|  8.92E-05|+/-1.04E-05|Jy|2005ApJS..161...41L|uncertainty|4.52       microns   | Broad-band measurement|171510.18 +600954.5 (J2000)| Flux in fixed aperture|Aperture =       7.59 arcsec.           |From new raw data
12|5.8 microns (IRAC)  | 74        |+/-19   | microJy            |5.23E+13|  7.40E-05|+/-1.90E-05|Jy|2007ApJ...664..713S|uncertainty|   5.731   microns   | Broad-band measurement|| Flux in fixed aperture|7.3" diameter aperture                  |From reprocessed raw data
13|5.8 microns (IRAC)  ||<100.00    |microJy             |5.23E+13||1.00E-04|Jy|2005ApJS..161...41L|3sigma plate limit|5.73       microns   | Broad-band measurement|171510.18 +600954.5 (J2000)| Flux in fixed aperture|Aperture =       7.59 arcsec.           |From new raw data
16|8.0 microns (IRAC)  | 149       |+/-27   | microJy            |3.81E+13|  1.49E-04|+/-2.70E-05|Jy|2007ApJ...664..713S|uncertainty|   7.872   microns   | Broad-band measurement|| Flux in fixed aperture|7.3" diameter aperture                  |From reprocessed raw data
17|8.0 microns (IRAC)  | 98.800    ||microJy             |3.81E+13|  9.88E-05||Jy|2007ApJ...658..778Y|no uncertainty reported|   7.872   microns   | Broad-band measurement|171510.28 +600955.2 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data
18|8.0 microns (IRAC)  | 153.12    |+/-21.29|microJy             |3.79E+13|  1.53E-04|+/-2.13E-05|Jy|2005ApJS..161...41L|uncertainty|7.91       microns   | Broad-band measurement|171510.18 +600954.5 (J2000)| Flux in fixed aperture|Aperture =       7.59 arcsec.           |From new raw data
19|8 microns (IRAC) | 2.8       |+/-1   %|milliJy             |3.75E+13|  2.80E-03|+/-2.80E-05|Jy|2009ApJ...698.1682W|typical accuracy|         8 microns   | Broad-band measurement|17 15 10.28 +60 09 55.2 (J2000)| Peak flux|                                        |From reprocessed raw data
1|MIPS 24um           | 1.50     |+/-0.45 |milliJy             |1.27E+13|  1.50E-03|+/-0.45E-03 |Jy|1996AJ....111.1431B|3sigma uncertainty|1.49       GHz       | Broad-band measurement| | Peak flux|                                        |From new raw data
21|24 microns (MIPS)   | 1.57      ||milliJy             |1.27E+13|  1.57E-03||Jy|2005ApJ...632L..13L|no uncertainty reported|   23.68   microns   | Broad-band measurement|17 15 10.28 +60 09 55.2 (J2000)| Total flux|                                        |From new raw data
22|24 microns (MIPS)   | 1500.852  ||microJy             |1.27E+13|  1.50E-03||Jy|2007ApJ...658..778Y|no uncertainty reported|   23.68   microns   | Broad-band measurement|171510.28 +600955.2 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data; measurementmodified from published value
2|MIPS 70um           | 5.0      |+/-1.4  |milliJy             |4.20E+12|  5.0E-03 |+/-1.4E-03|Jy|2010Natur.464..733S|3sigma uncertainty|     71.42 microns   | Broad-band measurement|21 35 11.6 -01 02 52.0 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
23|70 microns (MIPS)   | 5.7       |+/-1.2  | milliJy            |4.20E+12|  5.70E-03|+/-1.20E-03|Jy|2007ApJ...664..713S|estimated error|   71.42   microns   | Broad-band measurement|| Flux in fixed aperture|3 pixel radius aperture                 |From reprocessed raw data
3|MIPS 160um          |          |<30     |milliJy             |1.92E+12|          |30.0E-03|Jy|2009A&A...502..541E|3 sigma|     155.9 microns   | Broad-band measurement| | Flux in fixed aperture|                                        |From reprocessed raw data
4|MAMBO 1200um        | 0.99     |+/-0.43 |milliJy             |2.50E+11|  0.99E-03|+/-0.43E-03|Jy|2004MNRAS.354..779G|3sigma uncertainty|      1200 microns   | Broad-band measurement|16 37 06.7 +40 53 15 (J2000)| Flux integrated from map|S/N = 3.81                              |From new raw data
5|VLA 1.4GHz          |          |<0.08   |milliJy             |1.4E9   |          |0.08E-3 |Jy |2003MNRAS.343..293M|3sigma uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
