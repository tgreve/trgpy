
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-06-16T17:18:24PDT



Photometric Data for [HB89] 2343+125:BX0513

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|G (WHT)             | 24.13     ||mag                 |6.38E+14|  8.09E-07||Jy|2006ApJ...647..128E|no uncertainty reported|    0.47   microns   | Broad-band measurement|| Flux in fixed aperture|                                        |Averaged from previously published data
2|[N II] 6549 (Keck)  ||<0.6E-17   |erg/s/cm^2^         |4.58E+14||6.00E+05|Jy-Hz|2009ApJ...697.2057L|3 sigma|      6549 A         | Line measurement; flux integrated over line; lines measured in emission|23 46 11.133 +12 48 32.54 (J2000)| Flux integrated from map|                                        |From new raw data
3|H{alpha} (Keck II)  | 10.1E-17  |+/-0.4E-17|erg s^-1^ cm^-2^    |4.57E+14|  1.01E+07|+/-4.00E+05|Jy-Hz|2006ApJ...646..107E|uncertainty|    6563   A         | Line measurement; flux integrated over line; lines measured in emission|23 46 11.13 +12 48 32.14 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
4|H{alpha} (Keck)     | 5.4E-17   |+/-0.2E-17|erg/s/cm^2^         |4.57E+14|  5.40E+06|+/-2.00E+05|Jy-Hz|2009ApJ...697.2057L|1 sigma|      6563 A         | Line measurement; flux integrated over line; lines measured in emission|23 46 11.133 +12 48 32.54 (J2000)| Flux integrated from map|                                        |From new raw data
5|H{alpha} (VLT)      | 12.5E-17  |+/-1.8E-17|erg/s/cm^2^         |4.57E+14|  1.25E+07|+/-1.80E+06|Jy-Hz|2009ApJ...706.1364F|uncertainty|      6563 A         | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|                                        |From new raw data
6|[N II] 6585 (Keck)  | 1.8E-17   |+/-0.2E-17|erg/s/cm^2^         |4.55E+14|  1.80E+06|+/-2.00E+05|Jy-Hz|2009ApJ...697.2057L|1 sigma|      6585 A         | Line measurement; flux integrated over line; lines measured in emission|23 46 11.133 +12 48 32.54 (J2000)| Flux integrated from map|                                        |From new raw data
7|J (Hale/WIRC)       | 21.97     ||mag                 |2.40E+14|  2.54E-06||Jy|2006ApJ...646..107E|no uncertainty reported|    1.25   microns   | Broad-band measurement|23 46 11.13 +12 48 32.14 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data; derived from aflux in a different band and a color
8|K_s (Hale/WIRC)     | 20.10     ||mag                 |1.39E+14|  6.11E-06||Jy|2006ApJ...646..107E|no uncertainty reported|    2.15   microns   | Broad-band measurement|23 46 11.13 +12 48 32.14 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data
