
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-03-28T11:12:56PDT



Photometric Data for FFN 228

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|4.0-8 keV (Chandra) | |<0.22E-15  |ergs cm^-2^ s^-1^   |1.45E+18| |1.52E-11|Jy|2003AJ....126..539A|3 sigma|       6   keV       | Broad-band measurement|12 36 34.50 +62 12 41.2 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
2|4-8 keV (Chandra)   | |<0.36E-15  |erg cm^-2^ s^-1^    |1.45E+18| |2.48E-11|Jy|2001AJ....122.2810B|no uncertainty reported|       6   keV       | Broad-band measurement|12 36 34.51 +62 12 41.6 (J2000)| Flux in fixed aperture|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
3|2-10 keV (Chandra)  | 1.74E-16  | |erg/cm^2^/s         |1.45E+18|  1.20E-11| |Jy|2010MNRAS.401.2763L|no uncertainty reported|      6.00 keV       | Broad-band measurement|189.143590 62.211280 (J2000)| Modelled datum|                                        |From reprocessed raw data; NED frequency assigned tomid-point of band in keV
4|2-8 keV (Chandra)   | |<0.27E-15  |erg cm^-2^ s^-1^    |1.21E+18| |2.23E-11|Jy|2001AJ....122.2810B|no uncertainty reported|       5   keV       | Broad-band measurement|12 36 34.51 +62 12 41.6 (J2000)| Flux in fixed aperture|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
5|2-8 keV (Chandra)   | |<17.4E-17  |erg/cm^2^/s         |1.21E+18| |1.44E-11|Jy|2009ApJ...698.1380M|no uncertainty reported|      5.00 keV       | Broad-band measurement|12 36 34.51 +62 12 40.9 (J2000)| Not reported in paper|                                        |Averaged from previously published data; NED frequencyassigned to mid-point of band in keV
6|2.0-8 keV (Chandra) | |<0.17E-15  |ergs cm^-2^ s^-1^   |1.21E+18| |1.41E-11|Jy|2003AJ....126..539A|3 sigma|       5   keV       | Broad-band measurement|12 36 34.50 +62 12 41.2 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
7|0.5-8 keV (Chandra) | 0.31E-15  |+/-4   %|erg cm^-2^ s^-1^    |1.03E+18|  3.01E-11|+/-1.20E-12|Jy|2001AJ....122.2810B|estimated error|    4.25   keV       | Broad-band measurement|12 36 34.51 +62 12 41.6 (J2000)| Flux in fixed aperture|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
8|0.5-8 keV (Chandra) | 28.9E-17  | |erg/cm^2^/s         |1.03E+18|  2.81E-11| |Jy|2009ApJ...698.1380M|no uncertainty reported|      4.25 keV       | Broad-band measurement|12 36 34.51 +62 12 40.9 (J2000)| Not reported in paper|                                        |Averaged from previously published data; NED frequencyassigned to mid-point of band in keV
9|0.5-8 keV (Chandra) | 0.29E-15  | |ergs cm^-2^ s^-1^   |1.03E+18|  2.82E-11| |Jy|2003AJ....126..539A|no uncertainty reported|    4.25   keV       | Broad-band measurement|12 36 34.50 +62 12 41.2 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
10|2.0-4 keV (Chandra) | 0.10E-15  | |ergs cm^-2^ s^-1^   |7.25E+17|  1.38E-11| |Jy|2003AJ....126..539A|no uncertainty reported|       3   keV       | Broad-band measurement|12 36 34.50 +62 12 41.2 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
11|1.0-2 keV (Chandra) | 0.06E-15  | |ergs cm^-2^ s^-1^   |3.63E+17|  1.65E-11| |Jy|2003AJ....126..539A|no uncertainty reported|     1.5   keV       | Broad-band measurement|12 36 34.50 +62 12 41.2 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
12|0.5-2 keV (Chandra) | 0.10E-15  | |ergs cm^-2^ s^-1^   |3.02E+17|  3.31E-11| |Jy|2003AJ....126..539A|no uncertainty reported|    1.25   keV       | Broad-band measurement|12 36 34.50 +62 12 41.2 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
13|0.5-2 keV (Chandra) | 0.10E-15  |+/-4   %|erg cm^-2^ s^-1^    |3.02E+17|  3.31E-11|+/-1.32E-12|Jy|2001AJ....122.2810B|estimated error|    1.25   keV       | Broad-band measurement|12 36 34.51 +62 12 41.6 (J2000)| Flux in fixed aperture|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
14|0.5-1 keV (Chandra) | 0.05E-15  | |ergs cm^-2^ s^-1^   |1.81E+17|  2.76E-11| |Jy|2003AJ....126..539A|no uncertainty reported|    0.75   keV       | Broad-band measurement|12 36 34.50 +62 12 41.2 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
15|U (KPNO) AB         | 24.3      | | mag                |8.22E+14|  6.92E-07| |Jy|2004AJ....127.3137C|no uncertainty reported| 3647.65   A         | Broad-band measurement|189.143890 +62.21148 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
16|B (Subaru) AB       | 24.1      | | mag                |6.77E+14|  8.32E-07| |Jy|2004AJ....127.3137C|no uncertainty reported| 4427.60   A         | Broad-band measurement|189.143890 +62.21148 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
17|V (Subaru) AB       | 23.9      | | mag                |5.48E+14|  1.00E-06| |Jy|2004AJ....127.3137C|no uncertainty reported| 5471.22   A         | Broad-band measurement|189.143890 +62.21148 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
18|R (Keck II) AB      | 23.70     | | mag                |4.62E+14|  1.20E-06| |Jy|2004AJ....127.3121W|no uncertainty reported|   648.7   A         | Broad-band measurement|12 36 34.540 +62 12 41.02 (J2000)| Total flux|                                        |From new raw data
19|R (Subaru) AB       | 23.4      | | mag                |4.59E+14|  1.59E-06| |Jy|2004AJ....127.3137C|no uncertainty reported| 6534.16   A         | Broad-band measurement|189.143890 +62.21148 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
20|R (SUBARU) AB       | 23.32     | |mag                 |4.58E+14|  1.71E-06| |Jy|2007MNRAS.377..203G|no uncertainty reported|    6550   A         | Broad-band measurement|12 36 34.50 +62 12 41.2 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
21|I (Cousins)         | 22.22     |+/-0.02 |mag                 |3.79E+14|  3.30E-06|+/-6.14E-08|Jy|2004ApJ...616...71S|1 sigma|    7900   A         | Broad-band measurement| | Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
22|I (Subaru) AB       | 22.7      | | mag                |3.76E+14|  3.02E-06| |Jy|2004AJ....127.3137C|no uncertainty reported| 7975.89   A         | Broad-band measurement|189.143890 +62.21148 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
23|z' (Subaru) AB      | 22.2      | | mag                |3.31E+14|  4.79E-06| |Jy|2004AJ....127.3137C|no uncertainty reported| 9069.21   A         | Broad-band measurement|189.143890 +62.21148 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
24|J (2MASS)           | 20.63     |+/-0.04 |mag                 |2.40E+14|  8.91E-06|+/-3.34E-07|Jy|2004ApJ...616...71S|1 sigma|    1.25   microns   | Broad-band measurement| | Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
25|HK' (UH) AB         | 20.8      | | mag                |1.58E+14|  1.74E-05| |Jy|2004AJ....127.3137C|no uncertainty reported|18947.38   A         | Broad-band measurement|189.143890 +62.21148 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
26|K_s_ (2MASS)        | 18.51     |+/-0.03 |mag                 |1.38E+14|  2.63E-05|+/-7.37E-07|Jy|2004ApJ...616...71S|1 sigma|    2.17   microns   | Broad-band measurement| | Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
27|3.6 microns (IRAC)  | 62.42     |+/-0.06 |microJy             |8.44E+13|  6.24E-05|+/-6.00E-08|Jy|2007MNRAS.377..203G|uncertainty|   3.550   microns   | Broad-band measurement|12 36 34.50 +62 12 41.2 (J2000)| Corrected to total flux from single aperture measurement|                                        |From reprocessed raw data
28|3.6 microns (IRAC)  | 66.2      |+/-6.8  |microJy             |8.44E+13|  6.62E-05|+/-6.80E-06|Jy|2009ApJ...699.1610H|uncertainty|     3.550 microns   | Broad-band measurement|12 36 34.54 +62 12 41.1 (J2000)| Flux in fixed aperture|                                        |From new raw data
29|3.6 microns (IRAC)  | 64.50     |+/-3.23 |microJy             |8.44E+13|  6.45E-05|+/-3.23E-06|Jy|2011AJ....141....1T|rms uncertainty|     3.550 microns   | Broad-band measurement|189.143799 62.211391 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
30|4.5 microns (IRAC)  | 71.51     |+/-0.08 |microJy             |6.67E+13|  7.15E-05|+/-8.00E-08|Jy|2007MNRAS.377..203G|uncertainty|   4.493   microns   | Broad-band measurement|12 36 34.50 +62 12 41.2 (J2000)| Corrected to total flux from single aperture measurement|                                        |From reprocessed raw data
31|4.5 microns (IRAC)  | 74.5      |+/-7.6  |microJy             |6.67E+13|  7.45E-05|+/-7.60E-06|Jy|2009ApJ...699.1610H|uncertainty|     4.493 microns   | Broad-band measurement|12 36 34.54 +62 12 41.1 (J2000)| Flux in fixed aperture|                                        |From new raw data
32|4.5 microns (IRAC)  | 71.30     |+/-3.57 |microJy             |6.67E+13|  7.13E-05|+/-3.57E-06|Jy|2011AJ....141....1T|rms uncertainty|     4.493 microns   | Broad-band measurement|189.143799 62.211391 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
33|5.8 microns (IRAC)  | 58.82     |+/-0.44 |microJy             |5.23E+13|  5.88E-05|+/-4.40E-07|Jy|2007MNRAS.377..203G|uncertainty|   5.731   microns   | Broad-band measurement|12 36 34.50 +62 12 41.2 (J2000)| Corrected to total flux from single aperture measurement|                                        |From reprocessed raw data
34|5.8 microns (IRAC)  | 60.8      |+/-6.2  |microJy             |5.23E+13|  6.08E-05|+/-6.20E-06|Jy|2009ApJ...699.1610H|uncertainty|     5.731 microns   | Broad-band measurement|12 36 34.54 +62 12 41.1 (J2000)| Flux in fixed aperture|                                        |From new raw data
35|5.8 microns (IRAC)  | 58.00     |+/-2.93 |microJy             |5.23E+13|  5.80E-05|+/-2.93E-06|Jy|2011AJ....141....1T|rms uncertainty|     5.731 microns   | Broad-band measurement|189.143799 62.211391 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
36|8.0 microns (IRAC)  | 75.7      |+/-7.8  |microJy             |3.85E+13|  7.57E-05|+/-7.80E-06|Jy|2009ApJ...699.1610H|uncertainty|     7.782 microns   | Broad-band measurement|12 36 34.54 +62 12 41.1 (J2000)| Flux in fixed aperture|                                        |From new raw data
37|8.0 microns (IRAC)  | 70.47     |+/-0.45 |microJy             |3.81E+13|  7.05E-05|+/-4.50E-07|Jy|2007MNRAS.377..203G|uncertainty|   7.872   microns   | Broad-band measurement|12 36 34.50 +62 12 41.2 (J2000)| Corrected to total flux from single aperture measurement|                                        |From reprocessed raw data
38|8.0 microns (IRAC)  | 70.50     |+/-3.55 |microJy             |3.81E+13|  7.05E-05|+/-3.55E-06|Jy|2011AJ....141....1T|rms uncertainty|     7.872 microns   | Broad-band measurement|189.143799 62.211391 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
39|11 microns (AKARI)  | 104.0     |+/-15   | microJy            |2.73E+13|  1.04E-04|+/-1.50E-05|Jy|2009MNRAS.394..375N|uncertainty|        11 microns   | Broad-band measurement|12 36 34.53 +62 12 41.34 (J2000)| Flux integrated from map|                                        |From new raw data
40|ISOCAM 15 microns   | 0.4442    |+/-0.1  |milliJy             |2.07E+13|  4.44E-04|+/-1.00E-04|Jy|1997MNRAS.289..465G|estimated error|14.5       microns   | Broad-band measurement|123634.37 +621238.6 (J2000)| Flux integrated from map|                                        |From new raw data
41|15 microns (ISOCAM) | 363       |+/-60   |microJy             |2.00E+13|  3.63E-04|+/-6.00E-05|Jy|2006A&A...451...57M|68% confidence|    15.0   microns   | Broad-band measurement|189.1438751 62.2114830 (J2000)| Flux integrated from map|                                        |Averaged from previously published data
42|16 microns (IRS)    | 922.6     |+/-23.1 |microJy             |1.90E+13|  9.23E-04|+/-2.31E-05|Jy|2011AJ....141....1T|rms uncertainty|      15.8 microns   | Broad-band measurement|189.143799 62.211391 (J2000)| From fitting to map|                                        |From new raw data
43|16 microns (Spitzer)| 0.992     |+/-0.012| milliJy            |1.87E+13|  9.92E-04|+/-1.20E-05|Jy|2008ApJ...675.1171P|uncertainty|        16 microns   | Broad-band measurement|12 36 34.51 +62 12 40.9 (J2000)| Flux integrated from map|                                        |Averaged from previously published data
44|16 microns (IRS)    | 923       |+/-32   | microJy            |1.87E+13|  9.23E-04|+/-3.20E-05|Jy|2009MNRAS.394..375N|uncertainty|        16 microns   | Broad-band measurement|12 36 34.53 +62 12 41.34 (J2000)| Flux integrated from map|                                        |Averaged from previously published data
45|16 microns (Spitzer)| 993.6     | |microJy             |1.87E+13|  9.94E-04| |Jy|2009ApJ...698.1380M|no uncertainty reported|        16 microns   | Broad-band measurement|12 36 34.51 +62 12 40.9 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
46|18 microns (AKARI)  | 705       |+/-32   | microJy            |1.67E+13|  7.05E-04|+/-3.20E-05|Jy|2009MNRAS.394..375N|uncertainty|        18 microns   | Broad-band measurement|12 36 34.53 +62 12 41.34 (J2000)| Flux integrated from map|                                        |From new raw data
47|24 microns (Spitzer)| 446       | |microJy             |1.27E+13|  4.46E-04| |Jy|2009ApJ...698.1380M|no uncertainty reported|     23.68 microns   | Broad-band measurement|12 36 34.51 +62 12 40.9 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
48|24 microns (MIPS)   | 446       |+/-5    |microJy             |1.27E+13|  4.46E-04|+/-5.00E-06|Jy|2006A&A...451...57M|68% confidence|   23.68   microns   | Broad-band measurement|189.1438751 62.2114830 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
49|24 microns (MIPS)   | 458.54    |+/-4.94 |microJy             |1.27E+13|  4.59E-04|+/-4.94E-06|Jy|2007MNRAS.377..203G|uncertainty|   23.68   microns   | Broad-band measurement|12 36 34.50 +62 12 41.2 (J2000)| Corrected to total flux from single aperture measurement|                                        |From reprocessed raw data
50|24 microns (MIPS)   | 442.0     |+/-46.0 |microJy             |1.27E+13|  4.42E-04|+/-4.60E-05|Jy|2009ApJ...699.1610H|uncertainty|     23.68 microns   | Broad-band measurement|123634.51 +621241.0 (J2000)| Flux in fixed aperture|                                        |From new raw data
51|24 microns (MIPS)   | 444.0     |+/-5.5  |microJy             |1.27E+13|  4.44E-04|+/-5.50E-06|Jy|2011AJ....141....1T|rms uncertainty|     23.68 microns   | Broad-band measurement|189.143799 62.211391 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
52|24 microns (Spitzer)| 446       |+/-5    |microJy             |1.27E+13|  4.46E-04|+/-5.00E-06|Jy|2011ApJ...726...93R|uncertainty|     23.68 microns   | Broad-band measurement|12 36 34.49 +62 12 41.0 (J2000)| Not reported in paper|                                        |Averaged from previously published data
53|24 microns (Spitzer)| 445       |+/-7    |microJy             |1.27E+13|  4.45E-04|+/-7.00E-06|Jy|2011ApJ...726...93R|uncertainty|     23.68 microns   | Broad-band measurement|12 36 34.49 +62 12 41.0 (J2000)| Not reported in paper|                                        |Averaged from previously published data
54|70 microns (Spitzer)| 13200     | |microJy             |4.20E+12|  1.32E-02| |Jy|2009ApJ...698.1380M|no uncertainty reported|     71.42 microns   | Broad-band measurement|12 36 34.51 +62 12 40.9 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
55|70 microns (Spitzer)| 13.9      |+/-1.8  | milliJy            |4.20E+12|  1.39E-02|+/-1.80E-03|Jy|2008ApJ...675.1171P|uncertainty|     71.42 microns   | Broad-band measurement|12 36 34.51 +62 12 40.9 (J2000)| Flux integrated from map|                                        |Averaged from previously published data
56|70 microns (MIPS)   | 13.9      |+/-1.8  |milliJy             |4.20E+12|  1.39E-02|+/-1.80E-03|Jy|2007ApJ...659..305H|uncertainty|   71.42   microns   | Broad-band measurement|12 36 34.51 +62 12 40.9 (J2000)| Flux integrated from map|Color corrected for galaxy SEDs         |From reprocessed raw data
57|70 microns (MIPS)   | 13.9      |+/-1.5  |milliJy             |4.20E+12|  1.39E-02|+/-1.50E-03|Jy|2009ApJ...699.1610H|uncertainty|     71.42 microns   | Broad-band measurement|123634.51 +621241.0 (J2000)| Flux in fixed aperture|                                        |From new raw data
58|70 microns (PACS)  | 13.2      |+/-0.7  |mJy                 |4.283E+12| 13.2E-03|+/-0.7E-03|Jy|2004MNRAS.354..779G|3sigma uncertainty|      1200 microns   | Broad-band measurement|16 36 55.9 +40 59 12 (J2000)| Flux integrated from map|S/N = 3.66                              |From new raw data
59|100 microns (PACS) | 34.2      |+/-0.6  |mJy                 |2.998e+12| 34.2E-03|+/-0.6E-03 |Jy|2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
60|160 microns (PACS) | 63.2      |+/-1.6  |mJy                 |1.874e+12| 63.2E-03 |+/-1.6E-03 |Jy|2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
61|160 microns (MIPS)  | 110       |+/-27   |milliJy             |1.92E+12|  1.10E-01|+/-2.70E-02|Jy|2007ApJ...659..305H|uncertainty|   155.9   microns   | Broad-band measurement|12 36 34.51 +62 12 40.9 (J2000)| Flux integrated from map|Color corrected for galaxy SEDs         |From reprocessed raw data
62|250 microns (SPIRE)| 62.5      |+/-3.7  |mJy                 |1.199e+12| 62.5E-03|+/-3.7e-03 |Jy|2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
63|350 microns (SPIRE)| 47.1      |+/-3.0  |mJy                 |8.565E+11| 47.1E-03|+/-3.0E-03|Jy|2004MNRAS.354..779G|3sigma uncertainty|      1200 microns   | Broad-band measurement|16 36 55.9 +40 59 12 (J2000)| Flux integrated from map|S/N = 3.66                              |From new raw data
64|500 microns (SPIRE)| 19.6      |+/-4.0  |mJy                 |5.996E+11| 19.6E-03|+/-4.0E-03|Jy|2004MNRAS.354..779G|3sigma uncertainty|      1200 microns   | Broad-band measurement|16 36 55.9 +40 59 12 (J2000)| Flux integrated from map|S/N = 3.66                              |From new raw data
65|850 microns (SCUBA) | 3.0       |+/-0.8  |milliJy             |3.53E+11|  3.00E-03|+/-8.00E-04|Jy|2005MNRAS.358..149P|uncertainty|     850   microns   | Broad-band measurement|12 36 35.5 +62 12 38 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
66|850 microns (SCUBA) | 2.2       |+/-0.8  |milliJy             |3.53E+11|  2.20E-03|+/-8.00E-04|Jy|2005MNRAS.358..149P|uncertainty|     850   microns   | Broad-band measurement|12 36 35.5 +62 12 38 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
67|850 microns (SCUBA) | 4.3       |+/-1.4  |milliJy             |3.53E+11|  4.30E-03|+/-1.40E-03|Jy|2005ApJ...622..772C|uncertainty|     850   microns   | Broad-band measurement|123634.51 +621241.0 (J2000)| Flux integrated from map|                                        |From new raw data
68|1160 microns (Penner)|         |<1.8    |mJy                 |2.58442E+11|       |1.8E-03|Jy|2004MNRAS.354..779G|3sigma uncertainty|      1200 microns   | Broad-band measurement|16 36 55.9 +40 59 12 (J2000)| Flux integrated from map|S/N = 3.66                              |From new raw data
69|8.5 GHz             | 38.50     | |microJy             |8.50E+09|  3.85E-05| |Jy|1998AJ....116.1039R|no uncertainty reported|8.5        GHz       | Broad-band measurement; peak value reported; synthetic band|123634.505 +621240.99 (J2000)| Flux integrated from map; Pointing and beam filling|                                        |From new raw data; Corrected for contaminating sources
70|8.5 GHz             | 38.50     | |microJy             |8.50E+09|  3.85E-05| |Jy|1998AJ....116.1039R|no uncertainty reported|8.5        GHz       | Broad-band measurement; broad-band flux derived by integration over spectrum; synthetic band|123634.505 +621240.99 (J2000)| Flux integrated from map; Pointing and beam filling|                                        |From new raw data; Corrected for contaminating sources
71|8.4 GHz             | 40        |+/-3    |uJy                 |8.40E+09|  4.00E-05|+/-3.00E-06|Jy|1997ApJ...475L...5F|estimated error| 8.4       GHz       | Broad-band measurement|123634.49 +621240.9 (J2000)| Flux integrated from map; Beam filling or dilution corrected|                                        |From new raw data
72|1.4 GHz (VLA)       | 178.62    | |microJy             |1.40E+09|  1.79E-04| |Jy|2006A&A...451...57M|no uncertainty reported|     1.4   GHz       | Broad-band measurement|189.1438751 62.2114830 (J2000)| Flux integrated from map|                                        |From new raw data
73|1.4 GHz (VLA)       | 201.1     |+/-10.3 |microJy             |1.40E+09|  2.01E-04|+/-1.03E-05|Jy|2010ApJS..188..178M|uncertainty|       1.4 GHz       | Broad-band measurement|12 36 34.49 +62 12 41.0 (J2000)| Total flux; Beam filling or dilution corrected|Major=0.8"; Minor=0.7"; PA=65 deg       |From new raw data
74|1.4 GHz (VLA)       | 188       |+/-12   | microJy            |1.40E+09|  1.88E-04|+/-1.20E-05|Jy|2006MNRAS.371..963B|1 sigma|       1.4 GHz       | Broad-band measurement|12 36 34.508 +62 12 41.00 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
75|1.4 GHz             | 230.0     |+/-13.8 |microJy             |1.40E+09|  2.30E-04|+/-1.38E-05|Jy|2000ApJ...533..611R|1 sigma|1.4        GHz       | Broad-band measurement; broad-band flux derived by integration over spectrum; synthetic band|123634.515 +621241.01 (J2000)| Flux integrated from map; Pointing and beam filling|                                        |From new raw data; Corrected for contaminating sources
76|1.4 GHz (VLA)       | 230       | |microJy             |1.40E+09|  2.30E-04| |Jy|2005MNRAS.358.1159M|no uncertainty reported|     1.4   GHz       | Broad-band measurement|12 36 34.5168 +62 12 41.107 (J2000)| Flux integrated from map|                                        |From new raw data
