
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-04-04T05:28:04PDT



Photometric Data for GOODS J123600.15+621047.5

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|2-8 keV (Chandra)   | |<34.1E-17  |erg/cm^2^/s         |1.21E+18| |2.82E-11|Jy|2009ApJ...698.1380M|no uncertainty reported|      5.00 keV       | Broad-band measurement|12 36 00.17 +62 10 47.3 (J2000)| Not reported in paper|                                        |Averaged from previously published data; NED frequencyassigned to mid-point of band in keV
2|0.5-8 keV (Chandra) | |<19.9E-17  |erg/cm^2^/s         |1.03E+18| |1.93E-11|Jy|2009ApJ...698.1380M|no uncertainty reported|      4.25 keV       | Broad-band measurement|12 36 00.17 +62 10 47.3 (J2000)| Not reported in paper|                                        |Averaged from previously published data; NED frequencyassigned to mid-point of band in keV
3|R (Keck II) AB      | 25.20     | | mag                |4.62E+14|  3.02E-07| |Jy|2004AJ....127.3121W|no uncertainty reported|   648.7   A         | Broad-band measurement|12 36 00.188 +62 10 47.35 (J2000)| Total flux|                                        |From new raw data
4|H{alpha} (Keck)     | 3.7E-19   |+/-0.3E-19| W/m^2^             |4.57E+14|  8.10E-08|+/-6.56E-09|Jy|2004ApJ...617...64S|uncertainty|      6563 A         | Line measurement; flux integrated over line; lines measured in emission|123600.15 +621047.2 (J2000)| Flux integrated from map|                                        |From new raw data
5|I (Cousins)         | 23.08     |+/-0.03 |mag                 |3.79E+14|  1.50E-06|+/-4.19E-08|Jy|2004ApJ...616...71S|1 sigma|    7900   A         | Broad-band measurement| | Flux in fixed aperture|4" aper; phot contam by near neighbor   |Averaged new and previously published data
6|J (2MASS)           | 21.17     |+/-0.10 |mag                 |2.40E+14|  5.42E-06|+/-5.23E-07|Jy|2004ApJ...616...71S|1 sigma|    1.25   microns   | Broad-band measurement| | Flux in fixed aperture|4" aper; phot contam by near neighbor   |Averaged new and previously published data
7|F160W (HST) AB      | 22.64     |+/-0.08 |mag                 |1.87E+14|  3.19E-06|+/-2.35E-07|Jy|2010MNRAS.405..234S|uncertainty|      1.60 microns   | Broad-band measurement|12 36 00.15 +62 10 47.2 (J2000)| Flux in fixed aperture|                                        |From new raw data
8|K_s_ (2MASS)        | 20.02     |+/-0.15 |mag                 |1.38E+14|  6.55E-06|+/-9.70E-07|Jy|2004ApJ...616...71S|1 sigma|    2.17   microns   | Broad-band measurement| | Flux in fixed aperture|4" aper; phot contam by near neighbor   |Averaged new and previously published data
9|3.6 microns (IRAC)  | 12.9      |+/-1.6  |microJy             |8.44E+13|  1.29E-05|+/-1.60E-06|Jy|2009ApJ...699.1610H|uncertainty|     3.550 microns   | Broad-band measurement|12 36 00.16 +62 10 47.3 (J2000)| Flux in fixed aperture|                                        |From new raw data
10|3.6 microns (IRAC)  | 12.90     |+/-0.65 |microJy             |8.44E+13|  1.29E-05|+/-6.50E-07|Jy|2011AJ....141....1T|rms uncertainty|     3.550 microns   | Broad-band measurement|189.000687 62.179832 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
11|4.5 microns (IRAC)  | 15.2      |+/-1.7  |microJy             |6.67E+13|  1.52E-05|+/-1.70E-06|Jy|2009ApJ...699.1610H|uncertainty|     4.493 microns   | Broad-band measurement|12 36 00.16 +62 10 47.3 (J2000)| Flux in fixed aperture|                                        |From new raw data
12|4.5 microns (IRAC)  | 14.80     |+/-0.74 |microJy             |6.67E+13|  1.48E-05|+/-7.40E-07|Jy|2011AJ....141....1T|rms uncertainty|     4.493 microns   | Broad-band measurement|189.000687 62.179832 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
13|5.8 microns (IRAC)  | 27.7      |+/-2.9  |microJy             |5.23E+13|  2.77E-05|+/-2.90E-06|Jy|2009ApJ...699.1610H|uncertainty|     5.731 microns   | Broad-band measurement|12 36 00.16 +62 10 47.3 (J2000)| Flux in fixed aperture|                                        |From new raw data
14|5.8 microns (IRAC)  | 26.70     |+/-1.41 |microJy             |5.23E+13|  2.67E-05|+/-1.41E-06|Jy|2011AJ....141....1T|rms uncertainty|     5.731 microns   | Broad-band measurement|189.000687 62.179832 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
15|8.0 microns (IRAC)  | 63.7      |+/-6.6  |microJy             |3.85E+13|  6.37E-05|+/-6.60E-06|Jy|2009ApJ...699.1610H|uncertainty|     7.782 microns   | Broad-band measurement|12 36 00.16 +62 10 47.3 (J2000)| Flux in fixed aperture|                                        |From new raw data
16|8.0 microns (IRAC)  | 59.10     |+/-3.00 |microJy             |3.81E+13|  5.91E-05|+/-3.00E-06|Jy|2011AJ....141....1T|rms uncertainty|     7.872 microns   | Broad-band measurement|189.000687 62.179832 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
17|16 microns (IRS)    | 461.3     |+/-23.7 |microJy             |1.90E+13|  4.61E-04|+/-2.37E-05|Jy|2011AJ....141....1T|rms uncertainty|      15.8 microns   | Broad-band measurement|189.000687 62.179832 (J2000)| From fitting to map|                                        |From new raw data
18|16 microns (Spitzer)| 0.478     |+/-0.011| milliJy            |1.87E+13|  4.78E-04|+/-1.10E-05|Jy|2008ApJ...675.1171P|uncertainty|        16 microns   | Broad-band measurement|12 36 00.16 +62 10 47.3 (J2000)| Flux integrated from map|                                        |Averaged from previously published data
19|16 microns (Spitzer)| 496.8     | |microJy             |1.87E+13|  4.97E-04| |Jy|2009ApJ...698.1380M|no uncertainty reported|        16 microns   | Broad-band measurement|12 36 00.17 +62 10 47.3 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
20|24 microns (Spitzer)| 1220      | |microJy             |1.27E+13|  1.22E-03| |Jy|2009ApJ...698.1380M|no uncertainty reported|     23.68 microns   | Broad-band measurement|12 36 00.17 +62 10 47.3 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
21|24 microns (MIPS)   | 1230.0    |+/-120.0|microJy             |1.27E+13|  1.23E-03|+/-1.20E-04|Jy|2009ApJ...699.1610H|uncertainty|     23.68 microns   | Broad-band measurement|123600.15 +621047.2 (J2000)| Flux in fixed aperture|                                        |From new raw data
22|24 microns (MIPS)   | 1144      | |microJy             |1.27E+13|  1.14E-03| |Jy|2010ApJ...719.1393D|no uncertainty reported|     23.68 microns   | Broad-band measurement|12 36 00.2 +62 10 47.3 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
23|24 microns (IRAC)   | 1237      |+/-8.0  | microJy            |1.27E+13|  1.24E-03|+/-8.00E-06|Jy|2009ApJ...691..560C|uncertainty|     23.68 microns   | Broad-band measurement|12 36 00.13 +62 10 47.2 (J2000)| Not reported in paper|                                        |Averaged from previously published data
24|24 microns (MIPS)   | 1240.0    |+/-10.2 |microJy             |1.27E+13|  1.24E-03|+/-1.02E-05|Jy|2011AJ....141....1T|rms uncertainty|     23.68 microns   | Broad-band measurement|189.000687 62.179832 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
25|70 microns (MIPS)   | |<3.8       |microJy             |4.20E+12| |3.80E-03|Jy|2009ApJ...699.1610H|3 sigma|     71.42 microns   | Broad-band measurement|123600.15 +621047.2 (J2000)| Flux in fixed aperture|                                        |From new raw data
26|70 microns (Spitzer)| 5.5       |+/-1.2  | milliJy            |4.20E+12|  5.50E-03|+/-1.20E-03|Jy|2008ApJ...675.1171P|uncertainty|     71.42 microns   | Broad-band measurement|12 36 00.16 +62 10 47.3 (J2000)| Flux integrated from map|                                        |Averaged from previously published data
27|70 microns (Spitzer)| 4030      | |milliJy             |4.20E+12|  4.03E-03| |Jy|2009ApJ...698.1380M|no uncertainty reported|     71.42 microns   | Broad-band measurement|12 36 00.17 +62 10 47.3 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
28|350 microns (SHARC2)| 22.3      |+/-6.3  |milliJy             |8.57E+11|  2.23E-02|+/-6.30E-03|Jy|2006ApJ...650..592K|uncertainty|     350   microns   | Broad-band measurement| | Total flux|                                        |From new raw data
29|850 microns (SCUBA) | 7.9       |+/-2.4  |milliJy             |3.53E+11|  7.90E-03|+/-2.40E-03|Jy|2005ApJ...622..772C|uncertainty|     850   microns   | Broad-band measurement|123600.15 +621047.2 (J2000)| Flux integrated from map|                                        |From new raw data
30|CO(3-2) line (IRAM) | |<1.3       |Jy km s^-1^         |3.46E+11| |4.86E-07|Jy|2005MNRAS.359.1165G|3 sigma|  1.9865             | Line measurement; flux integrated over line; lines measured in emission|... ... (J2000)| Flux integrated from map|                                        |From new raw data
31|1.4 GHz             | 131.0     |+/-10.6 |microJy             |1.40E+09|  1.31E-04|+/-1.06E-05|Jy|2000ApJ...533..611R|1 sigma|1.4        GHz       | Broad-band measurement; broad-band flux derived by integration over spectrum; synthetic band|123600.150 +621047.17 (J2000)| Flux integrated from map; Pointing and beam filling|                                        |From new raw data; Corrected for contaminating sources
32|1.4 GHz (VLA)       | 128.5     |+/-8.1  | microJy            |1.40E+09|  1.29E-04|+/-8.10E-06|Jy|2009ApJ...691..560C|uncertainty|       1.4 GHz       | Broad-band measurement|12 36 00.13 +62 10 47.2 (J2000)| Not reported in paper|                                        |From reprocessed raw data
33|1.4 GHz (VLA)       | 130.3     |+/-6.3  |microJy             |1.40E+09|  1.30E-04|+/-6.30E-06|Jy|2010ApJS..188..178M|uncertainty|       1.4 GHz       | Broad-band measurement|12 36 00.13 +62 10 47.2 (J2000)| Total flux; Beam filling or dilution corrected|Major=0.0"; Minor=0.0"; PA=0 deg        |From new raw data
34|1.4 GHz (VLA)       | 144       |+/-8    | microJy            |1.40E+09|  1.44E-04|+/-8.00E-06|Jy|2006MNRAS.371..963B|1 sigma|       1.4 GHz       | Broad-band measurement|12 36 00.142 +62 10 47.19 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
