

Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.


queryDateTime:2009-11-03T15:07:35PST






Photometric Data for MIPS8327 (z=2.441)

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|R (KPNO)            | 1.447     ||microJy             |4.66E+14|  1.45E-06||Jy|2007ApJ...658..778Y|no uncertainty reported|    6440   A         | Broad-band measurement|171535.78 +602825.5 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data
2|R (Cousins) m_aper  | 23.30     |+/-0.05 |mag                 |4.65E+14|  1.46E-06|+/-6.74E-08|Jy|2004AJ....128....1F|based on count statistics only|6440       A         | Broad-band measurement|171535.783 +602825.78 (J2000)| Flux in fixed aperture|3-arcsecond aperture                    |From new raw data
3|R (Cousins) m_aper  | 23.49     |+/-0.11 |mag                 |4.65E+14|  1.23E-06|+/-1.25E-07|Jy|2004AJ....128....1F|based on count statistics only|6440       A         | Broad-band measurement|171535.783 +602825.89 (J2000)| Flux in fixed aperture|3-arcsecond aperture                    |From new raw data
4|R (Cousins) m_tot   | 23.27     |+/-0.06 |mag                 |4.65E+14|  1.51E-06|+/-8.32E-08|Jy|2004AJ....128....1F|based on count statistics only|6440       A         | Broad-band measurement|171535.783 +602825.78 (J2000)| Total flux|                                        |From new raw data
5|R (Cousins) m_tot   | 23.42     |+/-0.11 |mag                 |4.65E+14|  1.31E-06|+/-1.33E-07|Jy|2004AJ....128....1F|based on count statistics only|6440       A         | Broad-band measurement|171535.783 +602825.89 (J2000)| Total flux|                                        |From new raw data
6|F160W (HST NICMOS)         | 20.95     ||mag                 |1.87E+14|  4.35E-06||Jy|2011ApJ...730..125Z|no uncertainty reported|      1.60 microns   | Broad-band measurement|| Flux integrated from map|                                        |From new raw data
7|F160W (HST NICMOS)         | 21.06     || mag                |1.86E+14|  3.93E-06||Jy|2008ApJ...680..232D|no uncertainty reported|      1.61 microns   | Broad-band measurement|17 15 35.62 +60 28 24.49 (J2000)| Flux integrated from map|                                        |From new raw data
8|3.6 microns (IRAC)  | 12        |+/-3    | microJy            |8.44E+13|  1.20E-05|+/-3.00E-06|Jy|2007ApJ...664..713S|uncertainty|   3.550   microns   | Broad-band measurement|| Flux in fixed aperture|7.3" diameter aperture                  |From reprocessed raw data
9|4.5 microns (IRAC)  | 7         |+/-4    | microJy            |6.67E+13|  7.00E-06|+/-4.00E-06|Jy|2007ApJ...664..713S|uncertainty|   4.493   microns   | Broad-band measurement|| Flux in fixed aperture|7.3" diameter aperture                  |From reprocessed raw data
13|8.0 microns (IRAC)  | 58.435    ||microJy             |3.81E+13|  5.84E-05||Jy|2007ApJ...658..778Y|no uncertainty reported|   7.872   microns   | Broad-band measurement|171535.78 +602825.5 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data
14|8.0 microns (IRAC)  | 46        |+/-25   | microJy            |3.81E+13|  4.60E-05|+/-2.50E-05|Jy|2007ApJ...664..713S|uncertainty|   7.872   microns   | Broad-band measurement|| Flux in fixed aperture|7.3" diameter aperture                  |From reprocessed raw data
15|8 microns (IRAC) | 1.5       |+/-1   %|milliJy             |3.75E+13|  1.50E-03|+/-1.50E-05|Jy|2009ApJ...698.1682W|typical accuracy|         8 microns   | Broad-band measurement|17 15 35.78 +60 28 25.5 (J2000)| Peak flux|                                        |From reprocessed raw data
16|24 microns (MIPS)   | 1144.055  ||microJy             |1.27E+13|  1.14E-03||Jy|2007ApJ...658..778Y|no uncertainty reported|   23.68   microns   | Broad-band measurement|171535.78 +602825.5 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data; measurementmodified from published value
1|MIPS 24um           | 1.16     |+/-0.35  |milliJy            |1.27E+13|  1.16E-03|+/-0.35E-03 |Jy|1996AJ....111.1431B|uncertainty|1.49       GHz       | Broad-band measurement| | Peak flux|                                        |From new raw data
2|MIPS 70um           |          |<5.8    |milliJy             |4.20E+12|          |5.8E-03|Jy|2010Natur.464..733S|3sigma uncertainty|     71.42 microns   | Broad-band measurement|21 35 11.6 -01 02 52.0 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
18|70 microns (MIPS)   | 5.5       |+/-1.9  | milliJy            |4.20E+12|  5.50E-03|+/-1.90E-03|Jy|2007ApJ...664..713S|estimated error|   71.42   microns   | Broad-band measurement|| Flux in fixed aperture|3 pixel radius aperture                 |From reprocessed raw data
3|MIPS 160um          |          |<30     |milliJy             |1.92E+12|          |30.0E-03|Jy|2009A&A...502..541E|3 sigma|     155.9 microns   | Broad-band measurement| | Flux in fixed aperture|                                        |From reprocessed raw data
4|MAMBO 1200um        | 1.03     |+/-0.59 |milliJy             |2.50E+11|  1.03E-03|+/-0.59E-03|Jy|2004MNRAS.354..779G|uncertainty|      1200 microns   | Broad-band measurement|16 37 06.7 +40 53 15 (J2000)| Flux integrated from map|S/N = 3.81                              |From new raw data
5|VLA 1.4GHz          | 1.4      |+/-0.06 |milliJy             |1.4E9   |  1.4E-03 |+/-0.06E-03|Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
6|GMRT 610MHz         | 3.44     |+/-0.14 |milliJy             |610.E6  |  3.44E-03|+/-0.14E-03 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
