
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-02-19T12:23:33PST

z=2.38530

Photometric Data for MM J163650+4057

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
8|I (Cousins)         | 21.83     |+/-0.02 |mag                 |3.79E+14|  4.73E-06|+/-8.79E-08|Jy|2004ApJ...616...71S|1 sigma|    7900   A         | Broad-band measurement| | Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
9|F160W (HST) AB (WFC) | 21.85     |+/-0.04 |mag                 |1.87E+14|  6.61E-06|+/-2.43E-07|Jy|2010MNRAS.405..234S|uncertainty|      1.60 microns   | Broad-band measurement|16 36 50.43 +40 57 34.5 (J2000)| Flux in fixed aperture|                                        |From new raw data
10|K_s_ (2MASS)        | 18.43     |+/-0.02 |mag                 |1.38E+14|  2.83E-05|+/-5.26E-07|Jy|2004ApJ...616...71S|1 sigma|    2.17   microns   | Broad-band measurement| | Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
11|K (GeminiN)         | 18.85     |+/-0.10 |mag                 |1.36E+14|  1.85E-05|+/-1.70E-06|Jy|2011MNRAS.412..295T|uncertainty|      2.21 microns   | Broad-band measurement|| Flux in fixed aperture|6" diameter aperture                    |From new raw data
11|3.6 microns (IRAC)  | 31.9      |+/-3.3  |microJy             |8.44E+13|  3.19E-05|+/-3.30E-06|Jy|2009ApJ...699.1610H|uncertainty|     3.550 microns   | Broad-band measurement|16 36 50.41 +40 57 34.3 (J2000)| Flux in fixed aperture|                                        |From new raw data
12|4.5 microns (IRAC)  | 37.9      |+/-3.9  |microJy             |6.67E+13|  3.79E-05|+/-3.90E-06|Jy|2009ApJ...699.1610H|uncertainty|     4.493 microns   | Broad-band measurement|16 36 50.41 +40 57 34.3 (J2000)| Flux in fixed aperture|                                        |From new raw data
13|5.8 microns (IRAC)  | 51.9      |+/-5.4  |microJy             |5.23E+13|  5.19E-05|+/-5.40E-06|Jy|2009ApJ...699.1610H|uncertainty|     5.731 microns   | Broad-band measurement|16 36 50.41 +40 57 34.3 (J2000)| Flux in fixed aperture|                                        |From new raw data
15|8.0 microns (IRAC)  | 66.8      |+/-6.8  |microJy             |3.85E+13|  6.68E-05|+/-6.80E-06|Jy|2009ApJ...699.1610H|uncertainty|     7.782 microns   | Broad-band measurement|16 36 50.41 +40 57 34.3 (J2000)| Flux in fixed aperture|                                        |From new raw data
16|24 microns (MIPS)   | 1.02      |+/-10  %|milliJy             |1.27E+13|  1.02E-03|+/-1.02E-04|Jy|2009A&A...502..541E|uncertainty|     23.68 microns   | Broad-band measurement| | Flux in fixed aperture|                                        |From reprocessed raw data
17|24 microns (MIPS)   | 851.0     |+/-94.0 |microJy             |1.27E+13|  8.51E-04|+/-9.40E-05|Jy|2009ApJ...699.1610H|uncertainty|     23.68 microns   | Broad-band measurement|163650.43 +405734.5 (J2000)| Flux in fixed aperture|                                        |From new raw data
27|24 microns (MIPS)   | 9.8239E+02|+/-4.7230E+01|microJy             |1.27E+13|  9.82E-04|+/-4.72E-05|Jy|2013SSTSLC4.2....0C|uncertainty|23.68      microns   | Broad-band measurement|| Modelled datum|PSF fit                                 |From new raw data
28|24 microns (MIPS)   | 9.4716E+02|+/-4.4008E+01|microJy             |1.27E+13|  9.47E-04|+/-4.40E-05|Jy|2013SSTSLC4.2....0C|uncertainty|23.68      microns   | Broad-band measurement|| Flux in fixed aperture|14.7" aperture                          |From new raw data
18|70 microns (MIPS)   | |<5.5       |milliJy             |4.20E+12| |5.50E-03|Jy|2009A&A...502..541E|3 sigma|     71.42 microns   | Broad-band measurement| | Flux in fixed aperture|                                        |From reprocessed raw data
19|70 microns (MIPS)   | |<9.1       |milliJy             |4.20E+12| |9.10E-03|Jy|2009ApJ...699.1610H|3 sigma|     71.42 microns   | Broad-band measurement|163650.43 +405734.5 (J2000)| Flux in fixed aperture|                                        |From new raw data
20|160 microns (MIPS)  | |<22        |milliJy             |1.92E+12| |2.20E-02|Jy|2009A&A...502..541E|3 sigma|     155.9 microns   | Broad-band measurement| | Flux in fixed aperture|                                        |From reprocessed raw data
21|350 microns (SHARC2)| 33.0      |+/-5.6  |milliJy             |8.57E+11|  3.30E-02|+/-5.60E-03|Jy|2006ApJ...650..592K|uncertainty|     350   microns   | Broad-band measurement| | Total flux|                                        |From new raw data
23|850 microns (SCUBA) | 8.2       |+/-1.7  |milliJy             |3.53E+11|  8.20E-03|+/-1.70E-03|Jy|2005ApJ...622..772C|uncertainty|     850   microns   | Broad-band measurement|163650.43 +405734.5 (J2000)| Flux integrated from map|                                        |From new raw data
24|850 microns (SCUBA) | 8.3       |+/-1.8  |mag                 |3.53E+11|  8.30E-03|+/-1.80E-03|Jy|2006MNRAS.370.1057S|uncertainty|     850   microns   | Broad-band measurement|16 36 50.04 +40 57 33.0 (J2000)| From fitting to map|S/N = 5.20                              |From reprocessed raw data
26|1200 microns (MAMBO)| 3.1       |+/-0.7  | milliJy            |2.50E+11|  3.10E-03|+/-7.00E-04|Jy|2004MNRAS.354..779G|uncertainty|      1200 microns   | Broad-band measurement|16 36 50.3 +40 57 36 (J2000)| Flux integrated from map|S/N = 4.42                              |From new raw data
27|239.097 GHz (PdBI)  | 3.7       |+/-0.2  |milliJy             |2.39097E+11|  3.70E-03|+/-2.00E-04|Jy|2006ApJ...640..228T|uncertainty|     1.3   mm        | Broad-band measurement| | Flux integrated from map|                                        |From new raw data
27|1.3 mm (PdBI)       | 2.6       |+/-0.5  |milliJy             |2.31E+11|  2.60E-03|+/-5.00E-04|Jy|2006ApJ...640..228T|uncertainty|     1.3   mm        | Broad-band measurement| | Flux integrated from map|                                        |From new raw data
27|145.395 GHz (PdBI)  |           |<0.8  |milliJy             |1.45e+11| |8.00E-04|Jy|2006ApJ...640..228T|3 sigma|     1.3   mm        | Broad-band measurement| | Flux integrated from map|                                        |From new raw data
28|1.4 GHz (VLA)       | 216       |+/-12   | microJy            |1.40E+09|  2.16E-04|+/-1.20E-05|Jy|2006MNRAS.371..963B|1 sigma|       1.4 GHz       | Broad-band measurement|16 36 50.425 +40 57 34.45 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
29|1.4 GHz (VLA)       | 242       |+/-11   | microJy            |1.40E+09|  2.42E-04|+/-1.10E-05|Jy|2006MNRAS.371..963B|1 sigma|       1.4 GHz       | Broad-band measurement|16 36 50.425 +40 57 34.45 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
