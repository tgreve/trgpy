
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-06-11T08:35:35PDT



Photometric Data for BzK17999 (z=1.414)

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|R (Keck II) AB      | 24.88     | | mag                |4.62E+14|  4.05E-07| |Jy|2004AJ....127.3121W|no uncertainty reported|   648.7   A         | Broad-band measurement|12 37 51.859 +62 15 19.79 (J2000)| Total flux|                                        |From new raw data
2|3.6 microns (IRAC)  | 32.60     |+/-1.63 |microJy             |8.44E+13|  3.26E-05|+/-1.63E-06|Jy|2011AJ....141....1T|rms uncertainty|     3.550 microns   | Broad-band measurement|189.465881 62.255608 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
3|4.5 microns (IRAC)  | 35.90     |+/-1.80 |microJy             |6.67E+13|  3.59E-05|+/-1.80E-06|Jy|2011AJ....141....1T|rms uncertainty|     4.493 microns   | Broad-band measurement|189.465881 62.255608 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
4|5.8 microns (IRAC)  | 32.10     |+/-1.66 |microJy             |5.23E+13|  3.21E-05|+/-1.66E-06|Jy|2011AJ....141....1T|rms uncertainty|     5.731 microns   | Broad-band measurement|189.465881 62.255608 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
5|8.0 microns (IRAC)  | 37.10     |+/-1.92 |microJy             |3.81E+13|  3.71E-05|+/-1.92E-06|Jy|2011AJ....141....1T|rms uncertainty|     7.872 microns   | Broad-band measurement|189.465881 62.255608 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
6|16 microns (IRS)    | 238.6     |+/-8.3  |microJy             |1.90E+13|  2.39E-04|+/-8.30E-06|Jy|2011AJ....141....1T|rms uncertainty|      15.8 microns   | Broad-band measurement|189.465881 62.255608 (J2000)| From fitting to map|                                        |From new raw data
7|24 microns (MIPS)   | 226.0     |+/-4.8  |microJy             |1.27E+13|  2.26E-04|+/-4.80E-06|Jy|2011AJ....141....1T|rms uncertainty|     23.68 microns   | Broad-band measurement|189.465881 62.255608 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
7|24 microns (MIPS)   | 229.0     |+/-8.0  |microJy             |1.27E+13|  2.29E-04|+/-8.00E-06|Jy|2011AJ....141....1T|rms uncertainty|     23.68 microns   | Broad-band measurement|189.465881 62.255608 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
8|24 microns (Spitzer)| 230       |+/-8.0  |microJy             |1.27E+13|  2.30E-04|+/-8.0E-06 |Jy|2011ApJ...726...93R|no uncertainty reported|     23.68 microns   | Broad-band measurement|12 37 51.82 +62 15 20.2 (J2000)| Not reported in paper|                                        |Averaged from previously published data
11|70 microns (PACS)  |           |<2.0    |mJy                 |4.283E+12|         |2.0E-03|Jy|2004MNRAS.354..779G|3sigma uncertainty|      1200 microns   | Broad-band measurement|16 36 55.9 +40 59 12 (J2000)| Flux integrated from map|S/N = 3.66                              |From new raw data
10|100 microns (PACS) | 4.1       |+/-0.5  |microJy             |2.998e+12| 4.1E-03 |+/-0.5E-03 |Jy|2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
11|160 microns (PACS) | 10.8      |+/-1.4  |microJy             |1.874e+12| 10.8E-03|+/-1.4E-03 |Jy|2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
12|250 microns (SPIRE)| 14.7      |+/-2.5  |mJy                 |1.199e+12| 14.7E-03|+/-2.5e-03 |Jy|2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
13|350 microns (SPIRE)| 11.2      |+/-3.0  |mJy                 |8.565e+11| 11.2E-03|+/-3.0e-03 |Jy|2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
16|500 microns (SPIRE)|           |<12.0   |mJy                 |5.996E+11|         |12.0E-03|Jy|2004MNRAS.354..779G|3sigma uncertainty|      1200 microns   | Broad-band measurement|16 36 55.9 +40 59 12 (J2000)| Flux integrated from map|S/N = 3.66                              |From new raw data
15|1160 microns (Penner)|         |<1.8    |mJy                 |2.58442E+11|       |1.8E-03|Jy|2004MNRAS.354..779G|3sigma uncertainty|      1200 microns   | Broad-band measurement|16 36 55.9 +40 59 12 (J2000)| Flux integrated from map|S/N = 3.66                              |From new raw data
16|1.4 GHz (VLA)      | 28.3      |+/-5.6  |microJy             |1.40E+09|  2.83E-05|+/-5.60E-06|Jy|2010ApJS..188..178M|uncertainty|       1.4 GHz       | Broad-band measurement|12 37 51.82 +62 15 20.1 (J2000)| Total flux; Beam filling or dilution corrected|Major=0.0"; Minor=0.0"; PA=0 deg        |From new raw data
