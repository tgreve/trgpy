
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-07-10T07:43:22PDT



Photometric Data for PSS J2322+1944

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
2|I (HST)             | 17.92     ||mag                 |3.68E+14|  1.64E-04||Jy|2011ApJ...738...96M|no uncertainty reported|     0.814 microns   | Broad-band measurement|| Not reported in paper|                                        |From reprocessed raw data
3|F160W (HST/NIC2)    | 18.99     ||mag                 |1.87E+14|  2.75E-05||Jy|2006ApJ...649..616P|no uncertainty reported|   1.606   microns   | Broad-band measurement|23 22 07.02 +19 44 23 (J2000)| From fitting to map|Quasar mag; extinction = 0.03           |From new raw data; Extinction-corrected for Milky Way
5|3.6 microns (IRAC)  | 2.7550E+02|+/-4.1486E-01|microJy             |8.44E+13|  2.75E-04|+/-4.15E-07|Jy|2013SSTSLC4.2....0C|uncertainty|3.55       microns   | Broad-band measurement|| Flux in fixed aperture|5.8" aperture                           |From new raw data
6|3.6 microns (IRAC)  | 2.5506E+02|+/-3.8540E-01|microJy             |8.44E+13|  2.55E-04|+/-3.85E-07|Jy|2013SSTSLC4.2....0C|uncertainty|3.55       microns   | Broad-band measurement|| Flux in fixed aperture|3.8" aperture                           |From new raw data
7|4.5 microns (IRAC)  | 2.3915E+02|+/-4.4308E-01|microJy             |6.67E+13|  2.39E-04|+/-4.43E-07|Jy|2013SSTSLC4.2....0C|uncertainty|4.493      microns   | Broad-band measurement|| Flux in fixed aperture|3.8" aperture                           |From new raw data
8|4.5 microns (IRAC)  | 2.6057E+02|+/-5.4619E-01|microJy             |6.67E+13|  2.61E-04|+/-5.46E-07|Jy|2013SSTSLC4.2....0C|uncertainty|4.493      microns   | Broad-band measurement|| Flux in fixed aperture|5.8" aperture                           |From new raw data
9|5.8 microns (IRAC)  | 2.7648E+02|+/-1.3134E+00|microJy             |5.23E+13|  2.76E-04|+/-1.31E-06|Jy|2013SSTSLC4.2....0C|uncertainty|5.731      microns   | Broad-band measurement|| Flux in fixed aperture|3.8" aperture                           |From new raw data
10|5.8 microns (IRAC)  | 2.9061E+02|+/-1.6001E+00|microJy             |5.23E+13|  2.91E-04|+/-1.60E-06|Jy|2013SSTSLC4.2....0C|uncertainty|5.731      microns   | Broad-band measurement|| Flux in fixed aperture|5.8" aperture                           |From new raw data
11|8.0 microns (IRAC)  | 4.5984E+02|+/-2.2569E+00|microJy             |3.81E+13|  4.60E-04|+/-2.26E-06|Jy|2013SSTSLC4.2....0C|uncertainty|7.872      microns   | Broad-band measurement|| Flux in fixed aperture|3.8" aperture                           |From new raw data
12|8.0 microns (IRAC)  | 4.7043E+02|+/-2.9084E+00|microJy             |3.81E+13|  4.70E-04|+/-2.91E-06|Jy|2013SSTSLC4.2....0C|uncertainty|7.872      microns   | Broad-band measurement|| Flux in fixed aperture|5.8" aperture                           |From new raw data
13|24 microns (MIPS)   | 2.6887E+03|+/-2.1188E+01|microJy             |1.27E+13|  2.69E-03|+/-2.12E-05|Jy|2013SSTSLC4.2....0C|uncertainty|23.68      microns   | Broad-band measurement|| Modelled datum|PSF fit                                 |From new raw data
14|24 microns (MIPS)   | 2.5467E+03|+/-1.7950E+01|microJy             |1.27E+13|  2.55E-03|+/-1.80E-05|Jy|2013SSTSLC4.2....0C|uncertainty|23.68      microns   | Broad-band measurement|| Flux in fixed aperture|14.7" aperture                          |From new raw data
5|350 microns SHARC II| 79        |+/-11   |milliJy             |8.57E+11|  7.90E-02|+/-1.10E-02|Jy|2006ApJ...642..694B|1 sigma|     350   microns   | Broad-band measurement|23 22 07.25 +19 44 22.08 (J2000)| Flux integrated from map|                                        |From new raw data
18|850 microns (SCUBA) | 22.5      |+/-2.5 |milliJy             |3.53E+11|  22.5E-03|+/-2.5E-03|Jy|2007MNRAS.376.1073Z|no uncertainty reported|     850   microns   | Broad-band measurement|14 01 04.7 +02 52 28 (J2000)| Flux integrated from map|S/N = 9.6                               |From reprocessed raw data
7|1.2 mm (MAMBO)      | 9.6       |+/-0.5  | milliJy            |2.50E+11|  9.60E-03|+/-5.00E-04|Jy|2001A&A...374..371O|1 sigma|       1.2 mm        | Broad-band measurement|23 22 07.2 +19 44 23.0 (J2000)| Flux integrated from map|                                        |From new raw data
