
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2017-01-19T06:53:43PST



Photometric Data for NGC 0253

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
6|FUV (GALEX) AB      | 11.47     |+/-0.01 | mag                |1.98E+15|  9.38E-02|+/-8.64E-04|Jy|2007ApJS..173..185G|uncertainty|      1516 A         | Broad-band measurement|00 47 33.1 -25 17 17.6 (J2000)| Total flux|                                        |From new raw data
7|1530 A (GALEX) AB   | 11.01     |+/-0.02 |mag                 |1.96E+15|  1.43E-01|+/-2.64E-03|Jy|2006ApJS..164...38I|typical accuracy|    1530   A         | Broad-band measurement|00 47 26.14 -25 16 43.64 (J2000)| Total flux|                                        |From new raw data; Extinction-corrected for Milky Way
8|FUV (GALEX) AB      | 11.15     |+/-0.05 |mag                 |1.95E+15|  1.26E-01|+/-5.80E-03|Jy|2011ApJS..192....6L|uncertainty|      1539 A         | Broad-band measurement|| Flux in fixed aperture|                                        |From new raw data; Extinction-corrected for Milky Way
9|FUV (GALEX) AB      | 11.4603   |+/-0.00185201|mag                 |1.95E+15|  9.46E-02|+/-1.61E-04|Jy|2012GMSC..C...0000S|uncertainty|1538.6     A         | Broad-band measurement|11.888196279650 -25.28790532009 (J2000)| Flux integrated from map|Kron flux in elliptical aperture        |From new raw data
10|FUV (GALEX) AB      | 21.7563   |+/-0.269553|mag                 |1.95E+15|  7.20E-06|+/-1.79E-06|Jy|2012GMSC..C...0000S|uncertainty|1538.6     A         | Broad-band measurement|11.888196279650 -25.28790532009 (J2000)| Flux in fixed aperture|Flux in 7.5 arcsec diameter aperture    |From new raw data
11|1550 A (OAO)        | 9.08      |+/-0.55 |mag                 |1.93E+15|  6.80E-02|+/-4.48E-02|Jy|1982ApJ...256....1C|rms noise|1550       A         | Broad-band measurement|| Flux in fixed aperture|Aperture 10.0 arcmin                    |From new raw data
12|1910 A (OAO)        | 9.66      |+/-0.05 |mag                 |1.57E+15|  6.05E-02|+/-2.85E-03|Jy|1982ApJ...256....1C|rms noise|1910       A         | Broad-band measurement|| Flux in fixed aperture|Aperture 10.0 arcmin                    |From new raw data
13|NUV (GALEX) AB      | 10.94     |+/-0.01 | mag                |1.32E+15|  1.53E-01|+/-1.41E-03|Jy|2007ApJS..173..185G|uncertainty|      2267 A         | Broad-band measurement|00 47 33.1 -25 17 17.6 (J2000)| Total flux|                                        |From new raw data
14|2315 A (GALEX) AB   | 10.44     |+/-0.01 |mag                 |1.30E+15|  2.42E-01|+/-2.23E-03|Jy|2006ApJS..164...38I|typical accuracy|    2315   A         | Broad-band measurement|00 47 26.14 -25 16 43.64 (J2000)| Total flux|                                        |From new raw data; Extinction-corrected for Milky Way
15|NUV (GALEX) AB      | 10.8263   |+/-0.00047376|mag                 |1.29E+15|  1.70E-01|+/-7.40E-05|Jy|2012GMSC..C...0000S|uncertainty|2315.7     A         | Broad-band measurement|11.888196279650 -25.28790532009 (J2000)| Flux integrated from map|Kron flux in elliptical aperture        |From new raw data
16|NUV (GALEX) AB      | 20.9177   |+/-0.0612547|mag                 |1.29E+15|  1.56E-05|+/-8.80E-07|Jy|2012GMSC..C...0000S|uncertainty|2315.7     A         | Broad-band measurement|11.888196279650 -25.28790532009 (J2000)| Flux in fixed aperture|Flux in 7.5 arcsec diameter aperture    |From new raw data
17|NUV (GALEX) AB      | 10.62     |+/-0.03 |mag                 |1.29E+15|  2.05E-01|+/-5.67E-03|Jy|2011ApJS..192....6L|uncertainty|      2316 A         | Broad-band measurement|| Flux in fixed aperture|                                        |From new raw data; Extinction-corrected for Milky Way
18|2460 A (OAO)        | 9.64      |+/-0.03 |mag                 |1.22E+15|  1.02E-01|+/-2.86E-03|Jy|1982ApJ...256....1C|rms noise|2460       A         | Broad-band measurement|| Flux in fixed aperture|Aperture 10.0 arcmin                    |From new raw data
19|2980 A (OAO)        | 9.26      |+/-0.08 |mag                 |1.01E+15|  2.13E-01|+/-1.63E-02|Jy|1982ApJ...256....1C|rms noise|2980       A         | Broad-band measurement|| Flux in fixed aperture|Aperture 10.0 arcmin                    |From new raw data
20|3320 A (OAO)        | 8.93      |+/-0.05 |mag                 |9.03E+14|  3.58E-01|+/-1.69E-02|Jy|1982ApJ...256....1C|rms noise|3320       A         | Broad-band measurement|| Flux in fixed aperture|Aperture 10.0 arcmin                    |From new raw data
21|4250 A (OAO)        | 8.10      |+/-0.03 |mag                 |7.05E+14|  1.26E+00|+/-3.53E-02|Jy|1982ApJ...256....1C|rms noise|4250       A         | Broad-band measurement|| Flux in fixed aperture|Aperture 10.0 arcmin                    |From new raw data
22|B (Cousins) (B_26)  | 8.19      |+/-0.09 |mag                 |6.81E+14|  2.25E+00|+/-1.94E-01|Jy|1989ESOLV.C...0000L|typical accuracy|4400       A         | Broad-band measurement; photometric system transformed|004507 -2533.9 (B1950)| Modelled datum|See ESO-LV catalog for warning flag.    |From new raw data
23|B (Cousins) (B_25)  | 8.23      |+/-0.09 |mag                 |6.81E+14|  2.17E+00|+/-1.88E-01|Jy|1989ESOLV.C...0000L|typical accuracy|4400       A         | Broad-band measurement; photometric system transformed|004507 -2533.9 (B1950)| Modelled datum|See ESO-LV catalog for warning flag.    |From new raw data
24|B (B_T)             | 8.04      |+/-0.05 |mag                 |6.81E+14|  2.59E+00|+/-1.22E-01|Jy|1991RC3.9.C...0000d|rms uncertainty|4400       A         | Broad-band measurement|004505.7 -253340 (B1950)| Multiple methods|                                        |Homogenized from new and previously published data; StandardJohnson UBVRI filters assumed
25|B (m_B)             | 8.27      |+/-0.21 |mag                 |6.81E+14|  2.10E+00|+/-4.47E-01|Jy|1991RC3.9.C...0000d|rms uncertainty|4400       A         | Broad-band measurement|004505.7 -253340 (B1950)| Multiple methods|                                        |Homogenized from new and previously published data; StandardJohnson UBVRI filters assumed
26|B (Cousins) (B_T)   | 8.18      |+/-0.09 |mag                 |6.81E+14|  2.28E+00|+/-1.97E-01|Jy|1989ESOLV.C...0000L|typical accuracy|4400       A         | Broad-band measurement; photometric system transformed|004507 -2533.9 (B1950)| Modelled datum|See ESO-LV catalog for warning flag.    |From new raw data
27|B (B_T^0)           | 7.09      ||mag                 |6.81E+14|  6.21E+00||Jy|1991RC3.9.C...0000d|no uncertainty reported|4400       A         | Broad-band measurement|004505.7 -253340 (B1950)| Multiple methods|                                        |Homogenized from new and previously published data;Extinction-corrected for internal and Milky Way andK-correction applied; Standard Johnson UBVRI filtersassumed
28|B_J                 | 8.5247    ||mag                 |6.41E+14|  1.54E+00||Jy|2005MNRAS.361...34D|no uncertainty reported|    4680   A         | Broad-band measurement|004732.7 -251729.7 (J2000)| Flux in fixed aperture|                                        |From new raw data
29|R (Cousins) (R_25)  | 6.70      |+/-0.09 |mag                 |4.68E+14|  6.46E+00|+/-5.59E-01|Jy|1989ESOLV.C...0000L|typical accuracy|6400       A         | Broad-band measurement; photometric system transformed|004507 -2533.9 (B1950)| Modelled datum|See ESO-LV catalog for warning flag.    |From new raw data
30|R (Cousins) (R_T)   | 6.66      |+/-0.09 |mag                 |4.68E+14|  6.71E+00|+/-5.80E-01|Jy|1989ESOLV.C...0000L|typical accuracy|6400       A         | Broad-band measurement; photometric system transformed|004507 -2533.9 (B1950)| Modelled datum|See ESO-LV catalog for warning flag.    |From new raw data
31|R (Cousins) (R_26)  | 6.66      |+/-0.09 |mag                 |4.68E+14|  6.65E+00|+/-5.74E-01|Jy|1989ESOLV.C...0000L|typical accuracy|6400       A         | Broad-band measurement; photometric system transformed|004507 -2533.9 (B1950)| Modelled datum|See ESO-LV catalog for warning flag.    |From new raw data
32|R                   | 7.9725    ||mag                 |4.68E+14|  1.99E+00||Jy|2005MNRAS.361...34D|no uncertainty reported|    6400   A         | Broad-band measurement|004732.7 -251729.7 (J2000)| Flux in fixed aperture|                                        |From new raw data
34|I (SSO)             | 5.53      |+/-0.07 |mag                 |3.88E+14|  1.57E+01|+/-1.01E+00|Jy|2011ApJ...733...75H|uncertainty|      7730 A         | Broad-band measurement|00 47 33.12 -25 17 17.6 (J2000)| Flux in fixed aperture|                                        |From new raw data
35|I                   | 8.0555    ||mag                 |3.79E+14|  1.53E+00||Jy|2005MNRAS.361...34D|no uncertainty reported|    7900   A         | Broad-band measurement|004732.7 -251729.7 (J2000)| Flux in fixed aperture|                                        |From new raw data
36|J (ESO/SPM)         | 320.8     |+/-21.36|milliJy             |2.50E+14|  3.21E-01|+/-2.14E-02|Jy|1995ApJ...453..616S|rms uncertainty|1.198      microns   | Broad-band measurement|004505.7 -253337 (B1950)| Flux in fixed aperture|15" aperture                            |From new raw data
37|J (RGO)             | 8.6       |+/-0.09 |mag                 |2.50E+14|  5.95E-01|+/-5.15E-02|Jy|1973MNRAS.164..155G|uncertainty|       1.2 microns   | Broad-band measurement|| Flux in fixed aperture|25.2" aperture                          |From new raw data
38|J (Johnson)         | 6.81      |+/-0.03 |mag                 |2.42E+14|  3.03E+00|+/-8.48E-02|Jy|1977HarvU.T00M....A|uncertainty|   1.24    microns   | Broad-band measurement|| Flux in fixed aperture|105" aperture                           |From new raw data; derived from a flux in a different bandand a color
39|J_20 (2MASS LGA)    | 4.874     |+/-0.015|mag                 |2.40E+14|  1.79E+01|+/-2.49E-01|Jy|2003AJ....125..525J|1 sigma uncert.| 1.25      microns   | Broad-band measurement|004733.13 -251719.7 (J2000)| Flux integrated from map|1260.4 x  302.5 arcsec integration area.|From new raw data; Corrected for contaminating sources
40|J_Kron (2MASS LGA)  | 4.875     |+/-0.015|mag                 |2.40E+14|  1.79E+01|+/-2.48E-01|Jy|2003AJ....125..525J|1 sigma uncert.| 1.25      microns   | Broad-band measurement|004733.13 -251719.7 (J2000)| Flux integrated from map|1257.2 x  301.7 arcsec integration area.|From new raw data; Corrected for contaminating sources
41|J_tot (2MASS LGA)   | 4.814     |+/-0.016|mag                 |2.40E+14|  1.89E+01|+/-2.81E-01|Jy|2003AJ....125..525J|1 sigma uncert.| 1.25      microns   | Broad-band measurement|004733.13 -251719.7 (J2000)| Total flux|                                        |From new raw data
42|J_14arcsec (2MASS)  | 9.308     |+/-0.015|mag                 |2.40E+14|  3.01E-01|+/-4.19E-03|Jy|20032MASX.C.......:|1 sigma uncert.| 1.25      microns   | Broad-band measurement|004733.13 -251719.7 (J2000)| Flux in fixed aperture|14.0 x 14.0 arcsec aperture             |From new raw data
43|H (ESO/SPM)         | 640.0     |+/-42.62|milliJy             |1.90E+14|  6.40E-01|+/-4.26E-02|Jy|1995ApJ...453..616S|rms uncertainty|1.580      microns   | Broad-band measurement|004505.7 -253337 (B1950)| Flux in fixed aperture|15" aperture                            |From new raw data
44|H (RGO)             | 7.59      |+/-0.08 |mag                 |1.83E+14|  9.48E-01|+/-7.25E-02|Jy|1973MNRAS.164..155G|uncertainty|      1.64 microns   | Broad-band measurement|| Flux in fixed aperture|25.2" aperture                          |From new raw data
45|H_20 (2MASS LGA)    | 4.143     |+/-0.015|mag                 |1.82E+14|  2.25E+01|+/-3.14E-01|Jy|2003AJ....125..525J|1 sigma uncert.| 1.65      microns   | Broad-band measurement|004733.13 -251719.7 (J2000)| Flux integrated from map|1260.4 x  302.5 arcsec integration area.|From new raw data; Corrected for contaminating sources
46|H_Kron (2MASS LGA)  | 4.143     |+/-0.015|mag                 |1.82E+14|  2.25E+01|+/-3.14E-01|Jy|2003AJ....125..525J|1 sigma uncert.| 1.65      microns   | Broad-band measurement|004733.13 -251719.7 (J2000)| Flux integrated from map|1257.2 x  301.7 arcsec integration area.|From new raw data; Corrected for contaminating sources
47|H_tot (2MASS LGA)   | 4.088     |+/-0.016|mag                 |1.82E+14|  2.37E+01|+/-3.52E-01|Jy|2003AJ....125..525J|1 sigma uncert.| 1.65      microns   | Broad-band measurement|004733.13 -251719.7 (J2000)| Total flux|                                        |From new raw data
48|H_14arcsec (2MASS)  | 8.162     |+/-0.015|mag                 |1.82E+14|  5.57E-01|+/-7.74E-03|Jy|20032MASX.C.......:|1 sigma uncert.| 1.65      microns   | Broad-band measurement|004733.13 -251719.7 (J2000)| Flux in fixed aperture|14.0 x 14.0 arcsec aperture             |From new raw data
49|H (Johnson)         | 5.87      |+/-0.03 |mag                 |1.82E+14|  4.82E+00|+/-1.35E-01|Jy|1977HarvU.T00M....A|uncertainty|   1.65    microns   | Broad-band measurement|| Flux in fixed aperture|105" aperture                           |From new raw data; derived from a flux in a different bandand a color
50|H (HCO)             | 4.75      |+/-0.03 |mag                 |1.82E+14|  1.27E+01|+/-3.56E-01|Jy|1980ApJ...237..655A|uncertainty|   1.65    microns   | Broad-band measurement|| Flux in fixed aperture|316.5" aperture                         |From new raw data
51|H (HCO)             | 5.11      |+/-0.03 |mag                 |1.82E+14|  9.13E+00|+/-2.56E-01|Jy|1980ApJ...237..655A|uncertainty|   1.65    microns   | Broad-band measurement|| Flux in fixed aperture|212.8" aperture                         |From new raw data
52|H (HCO)             | 4.56      |+/-0.03 |mag                 |1.82E+14|  1.52E+01|+/-4.24E-01|Jy|1980ApJ...237..655A|uncertainty|   1.65    microns   | Broad-band measurement|| Flux in fixed aperture|409.6" aperture                         |From new raw data
53|1.65 microns        | 0.18      |+/-10  %|Jy                  |1.82E+14|  1.80E-01|+/-1.80E-02|Jy|1975ApJ...197...17R|uncertainty|    1.65   microns   | Broad-band measurement|| Flux in fixed aperture|5.5" aperture                           |From new raw data
56|K_20 (2MASS LGA)    | 3.822     |+/-0.016|mag                 |1.38E+14|  1.97E+01|+/-2.93E-01|Jy|2003AJ....125..525J|1 sigma uncert.| 2.17      microns   | Broad-band measurement|004733.13 -251719.7 (J2000)| Flux integrated from map|1260.4 x  302.5 arcsec integration area.|From new raw data; Corrected for contaminating sources
57|K_Kron (2MASS LGA)  | 3.823     |+/-0.016|mag                 |1.38E+14|  1.97E+01|+/-2.93E-01|Jy|2003AJ....125..525J|1 sigma uncert.| 2.17      microns   | Broad-band measurement|004733.13 -251719.7 (J2000)| Flux integrated from map|1257.2 x  301.7 arcsec integration area.|From new raw data; Corrected for contaminating sources
58|K_tot (2MASS LGA)   | 3.772     |+/-0.017|mag                 |1.38E+14|  2.07E+01|+/-3.26E-01|Jy|2003AJ....125..525J|1 sigma uncert.| 2.17      microns   | Broad-band measurement|004733.13 -251719.7 (J2000)| Total flux|                                        |From new raw data
59|K_s_14arcsec (2MASS)| 7.478     |+/-0.015|mag                 |1.38E+14|  6.80E-01|+/-9.47E-03|Jy|20032MASX.C.......:|1 sigma uncert.| 2.17      microns   | Broad-band measurement|004733.13 -251719.7 (J2000)| Flux in fixed aperture|14.0 x 14.0 arcsec aperture             |From new raw data
60|K (RGO)             | 6.9       |+/-0.07 |mag                 |1.37E+14|  1.13E+00|+/-7.52E-02|Jy|1973MNRAS.164..155G|uncertainty|      2.19 microns   | Broad-band measurement|| Flux in fixed aperture|25.2" aperture                          |From new raw data
61|2.2 microns         | 0.23      |+/-10  %|Jy                  |1.36E+14|  2.30E-01|+/-2.30E-02|Jy|1975ApJ...197...17R|uncertainty|     2.2   microns   | Broad-band measurement|| Flux in fixed aperture|5.5" aperture                           |From new raw data
62|K (ESO/SPM)         | 659.4     |+/-43.91|milliJy             |1.36E+14|  6.59E-01|+/-4.39E-02|Jy|1995ApJ...453..616S|rms uncertainty|2.210      microns   | Broad-band measurement|004505.7 -253337 (B1950)| Flux in fixed aperture|15" aperture                            |From new raw data
63|K (VLT)             | 12.34     ||mag                 |1.36E+14|  7.85E-03||Jy|2010ApJ...716.1166M|no uncertainty reported|     2.20  microns   | Broad-band measurement|| Flux in fixed aperture|Nucleus flux; 0.5" aperture             |From new raw data
64|K (Johnson)         | 5.46      |+/-0.03 |mag                 |1.35E+14|  4.37E+00|+/-1.22E-01|Jy|1977HarvU.T00M....A|uncertainty|   2.22    microns   | Broad-band measurement|| Flux in fixed aperture|105" aperture                           |From new raw data
65|L (RGO)             | 6.07      |+/-0.13 |mag                 |8.57E+13|  1.05E+00|+/-1.33E-01|Jy|1973MNRAS.164..155G|uncertainty|       3.5 microns   | Broad-band measurement|| Flux in fixed aperture|25.2" aperture                          |From new raw data
66|3.6 microns (IRAC)  | 1.26E+1   |+/-0.17E+1|Jy                  |8.44E+13|  1.26E+01|+/-1.70E+00|Jy|2009ApJ...703..517D|uncertainty|     3.550 microns   | Broad-band measurement|| Flux in fixed aperture|                                        |From reprocessed raw data; Extinction-corrected for Milky Way
67|3.6 microns         | 0.34      |+/-0.04 |Jy                  |8.33E+13|  3.40E-01|+/-4.00E-02|Jy|1975ApJ...197...17R|uncertainty|     3.6   microns   | Broad-band measurement|| Flux in fixed aperture|5.5" aperture                           |From new raw data
68|L (ESO/SPM)         | 858.4     |+/-57.17|milliJy             |7.95E+13|  8.58E-01|+/-5.72E-02|Jy|1995ApJ...453..616S|rms uncertainty|3.770      microns   | Broad-band measurement|004505.7 -253337 (B1950)| Flux in fixed aperture|15" aperture                            |From new raw data
69|4.5 microns (IRAC)  | 8.72E+0   |+/-1.20E+0|Jy                  |6.67E+13|  8.72E+00|+/-1.20E+00|Jy|2009ApJ...703..517D|uncertainty|     4.493 microns   | Broad-band measurement|| Flux in fixed aperture|                                        |From reprocessed raw data; Extinction-corrected for Milky Way
70|5.0 microns         | 3.2       |+/-1.1  |Jy                  |6.00E+13|  3.20E+00|+/-1.10E+00|Jy|1975ApJ...197...17R|uncertainty|     5.0   microns   | Broad-band measurement|| Flux in fixed aperture|13.5" aperture;Low quality data         |From new raw data
71|5.0 microns         | 0.37      |+/-0.06 |Jy                  |6.00E+13|  3.70E-01|+/-6.00E-02|Jy|1975ApJ...197...17R|uncertainty|     5.0   microns   | Broad-band measurement|| Flux in fixed aperture|5.5" aperture                           |From new raw data
72|5.8 microns (IRAC)  | 1.96E+1   |+/-0.24E+1|Jy                  |5.23E+13|  1.96E+01|+/-2.40E+00|Jy|2009ApJ...703..517D|uncertainty|     5.731 microns   | Broad-band measurement|| Flux in fixed aperture|                                        |From reprocessed raw data; Extinction-corrected for Milky Way
73|8.0 microns (IRAC)  | 4.54E+1   |+/-0.57E+1|Jy                  |3.81E+13|  4.54E+01|+/-5.70E+00|Jy|2009ApJ...703..517D|uncertainty|     7.872 microns   | Broad-band measurement|| Flux in fixed aperture|                                        |From reprocessed raw data; Extinction-corrected for Milky Way
74|8.8 microns         | 3         |+/-10  %|Jy                  |3.41E+13|  3.00E+00|+/-3.00E-01|Jy|1975ApJ...197...17R|uncertainty|     8.8   microns   | Broad-band measurement|| Flux in fixed aperture|5.5" aperture                           |From new raw data
75|8.9 microns TIMMI2  | 1140      |+/-15  %|milliJy             |3.37E+13|  1.14E+00|+/-1.71E-01|Jy|2008A&A...484..341R|estimated error|       8.9 microns   | Broad-band measurement|00 47 33.1 -25 17 17.2 (J2000)| Flux in fixed aperture|                                        |From new raw data
77|10 microns          | 6.20      |+/-0.3  |Jy                  |3.00E+13|  6.20E+00|+/-3.00E-01|Jy|1978ApJ...220L..37R|uncertainty|   10      microns   | Broad-band measurement|| Flux in fixed aperture|5.7" aperture                           |From new raw data
78|10 microns (IRTF)   | 6800      ||milliJy             |2.97E+13|  6.80E+00||Jy|1989ApJ...344..135H|no uncertainty reported|    10.1   microns   | Broad-band measurement|| Flux in fixed aperture|4" beam                                 |From new raw data
79|10.3 microns        | 2.9       |+/-10  %|Jy                  |2.91E+13|  2.90E+00|+/-2.90E-01|Jy|1975ApJ...197...17R|uncertainty|    10.3   microns   | Broad-band measurement|| Flux in fixed aperture|5.5" aperture                           |From new raw data
80|10.5 microns        | 6.2       |+/-0.5  |Jy                  |2.86E+13|  6.20E+00|+/-5.00E-01|Jy|1972ApJ...176L..95R|1 sigma|      10.5 microns   | Broad-band measurement|| Flux in fixed aperture|6" aperture                             |From new raw data
81|10.6 microns        | 6         |+/-10  %|Jy                  |2.83E+13|  6.00E+00|+/-6.00E-01|Jy|1975ApJ...197...17R|uncertainty|    10.6   microns   | Broad-band measurement|| Flux in fixed aperture|5.5" aperture                           |From new raw data
82|10.6 microns        | 10.5      |+/-10  %|Jy                  |2.83E+13|  1.05E+01|+/-1.05E+00|Jy|1975ApJ...197...17R|uncertainty|    10.6   microns   | Broad-band measurement|| Flux in fixed aperture|13.5" aperture                          |From new raw data
84|11.3 microns (IRS)  | 228E-20   |+/-68E-20| W/cm^2^            |2.65E+13|  2.28E+12|+/-6.80E+11|Jy-Hz|2004ApJS..154..242D|uncertainty|      11.3 microns   | Line measurement; flux integrated over line; lines measured in emission|00 47 33.2 -25 17 19 (J2000)| From fitting to map|Nuclear flux                            |From new raw data
85|11.6 microns        | 6.6       |+/-10  %|Jy                  |2.58E+13|  6.60E+00|+/-6.60E-01|Jy|1975ApJ...197...17R|uncertainty|    11.6   microns   | Broad-band measurement|| Flux in fixed aperture|5.5" aperture                           |From new raw data
87|12 microns (IRAS)   | 41.04     |+/-0.035|Jy                  |2.50E+13|  4.10E+01|+/-3.50E-02|Jy|2003AJ....126.1607S|1 sigma|      12   microns   | Broad-band measurement|00 47 33.1 -25 17 15 (J2000)| Total flux|Size, Method, Flag codes: RZ;see paper  |From reprocessed raw data
88|12.0 microns (IRS)  | 20E-20    |+/-6E-20| W/cm^2^            |2.50E+13|  2.00E+11|+/-6.00E+10|Jy-Hz|2004ApJS..154..242D|uncertainty|      12.0 microns   | Line measurement; flux integrated over line; lines measured in emission|00 47 33.2 -25 17 19 (J2000)| From fitting to map|Nuclear flux                            |From new raw data
89|12 microns (IRAS)   | 36.58     |+/-0.078|Jy                  |2.50E+13|  3.66E+01|+/-7.80E-02|Jy|1989AJ.....98..766S|rms noise|12         microns   | Broad-band measurement|004505.0 -253347 (B1950)| Integrated from scans|Resolved with 0.77' beam                |From reprocessed raw data
90|12 microns (IRAS)   | 2.402E+01 |+/-5   %|Jy                  |2.50E+13|  2.40E+01|+/-1.20E+00|Jy|1990IRASF.C...0000M|uncertainty| 12        microns   | Broad-band measurement|004505.7 -253337 (B1950)| Flux in fixed aperture|IRAS quality flag = 3                   |From new raw data
91|12 microns (IRAS)   | 55.84     |+/-25  %|Jy                  |2.50E+13|  5.58E+01|+/-1.40E+01|Jy|1988ApJS...68...91R|uncertainty|      12   microns   | Broad-band measurement|| Flux integrated from map|                                        |From reprocessed raw data
93|12.6 microns        | 11.2      |+/-10  %|Jy                  |2.38E+13|  1.12E+01|+/-1.12E+00|Jy|1975ApJ...197...17R|uncertainty|    12.6   microns   | Broad-band measurement|| Flux in fixed aperture|5.5" aperture                           |From new raw data
109|17 microns          | 23.5      |+/-6    |Jy                  |1.76E+13|  2.35E+01|+/-6.00E+00|Jy|1975ApJ...197...17R|uncertainty|      17   microns   | Broad-band measurement|| Flux in fixed aperture|5.5" aperture                           |From new raw data
115|19 microns          | 28        |+/-5    |Jy                  |1.58E+13|  2.80E+01|+/-5.00E+00|Jy|1975ApJ...197...17R|uncertainty|      19   microns   | Broad-band measurement|| Flux in fixed aperture|5.5" aperture                           |From new raw data
116|21 microns          | 56        |+/-20   |Jy                  |1.43E+13|  5.60E+01|+/-2.00E+01|Jy|1975ApJ...197...17R|uncertainty|      21   microns   | Broad-band measurement|| Flux in fixed aperture|13.5" aperture                          |From new raw data
117|21 microns          | 27        |+/-10  %|Jy                  |1.43E+13|  2.70E+01|+/-2.70E+00|Jy|1975ApJ...197...17R|uncertainty|      21   microns   | Broad-band measurement|| Flux in fixed aperture|5.5" aperture                           |From new raw data
118|22.5 microns        | 34        |+/-10  %|Jy                  |1.33E+13|  3.40E+01|+/-3.40E+00|Jy|1975ApJ...197...17R|uncertainty|    22.5   microns   | Broad-band measurement|| Flux in fixed aperture|5.5" aperture                           |From new raw data
119|24 microns (MIPS)   | 1.46E+2   |+/-0.16E+2|Jy                  |1.27E+13|  1.46E+02|+/-1.60E+01|Jy|2009ApJ...703..517D|uncertainty|     23.68 microns   | Broad-band measurement|| Flux in fixed aperture|                                        |From reprocessed raw data; Extinction-corrected for Milky Way
120|24 microns (MIPS)   | 140       ||Jy                  |1.27E+13|  1.40E+02||Jy|2005ApJ...628L..29E|no uncertainty reported|   23.68   microns   | Broad-band measurement|| Flux integrated from map|                                        |Transformed from previously published data
122|24.5 microns        | 52        |+/-10   |Jy                  |1.22E+13|  5.20E+01|+/-5.20E+00|Jy|1975ApJ...197...17R|uncertainty|    24.5   microns   | Broad-band measurement|| Flux in fixed aperture|5.5" aperture                           |From new raw data
123|25 microns (IRAS)   | 154.67    |+/-0.045|Jy                  |1.20E+13|  1.55E+02|+/-4.50E-02|Jy|2003AJ....126.1607S|1 sigma|      25   microns   | Broad-band measurement|00 47 33.1 -25 17 15 (J2000)| Total flux|Size, Method, Flag codes: RZ;see paper  |From reprocessed raw data
124|25 microns (IRAS)   | 137.89    |+/-0.194|Jy                  |1.20E+13|  1.38E+02|+/-1.94E-01|Jy|1989AJ.....98..766S|rms noise|25         microns   | Broad-band measurement|004505.0 -253347 (B1950)| Integrated from scans|Resolved with 0.78' beam                |From reprocessed raw data
125|25 microns (IRAS)   | 1.197E+02 |+/-7   %|Jy                  |1.20E+13|  1.20E+02|+/-1.68E+00|Jy|1990IRASF.C...0000M|uncertainty| 25        microns   | Broad-band measurement|004505.7 -253337 (B1950)| Flux in fixed aperture|IRAS quality flag = 3                   |From new raw data
126|25 microns (IRAS)   | 155.65    |+/-25  %|Jy                  |1.20E+13|  1.56E+02|+/-3.89E+01|Jy|1988ApJS...68...91R|uncertainty|      25   microns   | Broad-band measurement|| Flux integrated from map|                                        |From reprocessed raw data
137|34 microns          ||<200       |Jy                  |8.82E+12||2.00E+02|Jy|1975ApJ...197...17R|3sigma uncertainty|      34   microns   | Broad-band measurement|| Flux in fixed aperture|5.5" aperture                           |From new raw data
141|60 microns (ISO)    | 1044.7    |+/-20  %|Jy                  |5.00E+12|  1.04E+03|+/-2.09E+02|Jy|2001A&A...375..566N|uncertainty|      60   microns   | Broad-band measurement|| Modelled datum|                                        |From new raw data
142|60 microns (IRAS)   | 967.81    |+/-0.065|Jy                  |5.00E+12|  9.68E+02|+/-6.50E-02|Jy|2003AJ....126.1607S|1 sigma|      60   microns   | Broad-band measurement|00 47 33.1 -25 17 15 (J2000)| Total flux|Size, Method, Flag codes: RI;see paper  |From reprocessed raw data
143|60 microns (IRAS)   | 931.69    |+/-0.47 |Jy                  |5.00E+12|  9.32E+02|+/-4.70E-01|Jy|1989AJ.....98..766S|rms noise|60         microns   | Broad-band measurement|004505.0 -253347 (B1950)| Integrated from scans|Resolved with 1.44' beam                |From reprocessed raw data
144|60 microns (IRAS)   | 7.842E+02 |+/-6   %|Jy                  |5.00E+12|  7.84E+02|+/-4.71E+01|Jy|1990IRASF.C...0000M|uncertainty| 60        microns   | Broad-band measurement|004505.7 -253337 (B1950)| Flux in fixed aperture|IRAS quality flag = 3                   |From new raw data
145|60 microns (IRAS)   | 998.73    |+/-25  %|Jy                  |5.00E+12|  9.99E+02|+/-2.50E+02|Jy|1988ApJS...68...91R|uncertainty|      60   microns   | Broad-band measurement|| Flux integrated from map|                                        |From reprocessed raw data
148|70 microns (MIPS)   | 1.41E+3   |+/-0.17E+3|Jy                  |4.20E+12|  1.41E+03|+/-1.70E+02|Jy|2009ApJ...703..517D|uncertainty|     71.42 microns   | Broad-band measurement|| Flux in fixed aperture|                                        |From reprocessed raw data; Extinction-corrected for Milky Way
151|90 microns (AKARI)  | 1200      |+/-240  |Jy                  |3.33E+12|  1.20E+03|+/-2.40E+02|Jy|2009ApJ...698L.125K|uncertainty|        90 microns   | Broad-band measurement|00 47 33.1 -25 17 17.5 (J2000)| Flux in fixed aperture|Center flux                             |From new raw data
152|100 microns (IRAS)  | 1288.15   |+/-0.644|Jy                  |3.00E+12|  1.29E+03|+/-6.44E-01|Jy|2003AJ....126.1607S|1 sigma|     100   microns   | Broad-band measurement|00 47 33.1 -25 17 15 (J2000)| Total flux|Size, Method, Flag codes: RI;see paper  |From reprocessed raw data
153|100 microns (IRAS)  | 9.931E+02 |+/-7   %|Jy                  |3.00E+12|  9.93E+02|+/-6.95E+01|Jy|1990IRASF.C...0000M|uncertainty| 100       microns   | Broad-band measurement|004505.7 -253337 (B1950)| Flux in fixed aperture|IRAS quality flag = 2                   |From new raw data
154|100 microns (IRAS)  | 1861.67   |+/-25  %|Jy                  |3.00E+12|  1.86E+03|+/-4.65E+02|Jy|1988ApJS...68...91R|uncertainty|     100   microns   | Broad-band measurement|| Flux integrated from map|                                        |From reprocessed raw data
156|140 microns (AKARI) | 1300      |+/-390  |Jy                  |2.14E+12|  1.30E+03|+/-3.90E+02|Jy|2009ApJ...698L.125K|uncertainty|       140 microns   | Broad-band measurement|00 47 33.1 -25 17 17.5 (J2000)| Flux in fixed aperture|Center flux                             |From new raw data
159|160 microns (MIPS)  | 1.87E+3   |+/-0.29E+3|Jy                  |1.92E+12|  1.87E+03|+/-2.90E+02|Jy|2009ApJ...703..517D|uncertainty|     155.9 microns   | Broad-band measurement|| Flux in fixed aperture|                                        |From reprocessed raw data; Extinction-corrected for Milky Way
162|350 microns         | 172       |+/-51   |Jy                  |8.57E+11|  1.72E+02|+/-5.10E+01|Jy|1973ApJ...183L..67R|internal error| 350       microns   | Broad-band measurement|| Flux in fixed aperture|Beam diameter 63 arcsec                 |From new raw data
163|540 microns         | 25        |+/-10   |Jy                  |5.55E+11|  2.50E+01|+/-1.00E+01|Jy|1977ApJ...216..698H|estimated error| 540       microns   | Broad-band measurement|| Flux in fixed aperture|Beam diameter 83 arcsec                 |From new raw data
170|870 microns (LABOCA)| 17.6      |+/-1.8  |Jy                  |3.45E+11|  1.76E+01|+/-1.80E+00|Jy|2008A&A...490...77W|uncertainty|       870 microns   | Broad-band measurement|| Total flux|                                        |From new raw data
171|1 mm                | 4.4       |+/-1.7  |Jy                  |3.00E+11|  4.40E+00|+/-1.70E+00|Jy|1984A&A...137..117C|rms uncertainty|1          A         | Broad-band measurement; peak value reported|| Flux in fixed aperture|half-power beam width 3.9'              |From new raw data
172|1.25 mm (SEST)      | 4400.0    |+/-1700.0|milliJy             |2.40E+11|  4.40E+00|+/-1.70E+00|Jy|1996MNRAS.283...85A|uncertainty|    1.25   mm        | Broad-band measurement|00 45 05.2 -25 33 40 (B1950)| Flux integrated from map|From 1984A&A...137..117C                |Averaged from previously published data; K-correction applied
173|1.3 mm (NRAO)       | 0.7       |+/-0.3  |Jy                  |2.31E+11|  7.00E-01|+/-3.00E-01|Jy|1987ApJ...318..645T|uncertainty|       1.3 mm        | Broad-band measurement|00457.8 -253342 (B1950)| Not reported in paper|Beam size = 33"                         |From new raw data
174|2.6 mm (NRO)        | 120       |+/-30   | milliJy            |1.15E+11|  1.20E-01|+/-3.00E-02|Jy|2004ApJ...611..835P|uncertainty|      2.6  mm        | Broad-band measurement|| Peak flux|                                        |From new raw data
176|W (WMAP)            | 0.9       |+/-0.2  | Jy                 |9.40E+10|  9.00E-01|+/-2.00E-01|Jy|2009ApJS..180..283W|uncertainty|        94 GHz       | Broad-band measurement|00 47 19 -25 14 00 (J2000)| Flux integrated from map|                                        |From new raw data
177|94 GHz (WMAP)       | 0.7       |+/-0.4  |Jy                  |9.40E+10|  7.00E-01|+/-4.00E-01|Jy|2009ApJ...694..222C|1 sigma|        94 GHz       | Broad-band measurement|00 47 25 -25 16 00 (J2000)| Flux integrated from map|                                        |From new raw data
178|94 GHz (WMAP)       | 0.9       |+/-0.20 |Jy                  |9.40E+10|  9.00E-01|+/-2.00E-01|Jy|2011ApJS..192...15G|uncertainty|        94 GHz       | Broad-band measurement|00 47 20 -25 13 (J2000)| Flux integrated from map|                                        |From new raw data
185|61 GHz (WMAP)       | 1.9       |+/-0.6  |Jy                  |6.10E+10|  1.90E+00|+/-6.00E-01|Jy|2003ApJS..148...97B|uncertainty|      61   GHz       | Broad-band measurement|004717.7 -251228 (J2000)| Flux integrated from map|                                        |From new raw data
186|61 GHz (WMAP)       | 0.7       |+/-0.2  |Jy                  |6.10E+10|  7.00E-01|+/-2.00E-01|Jy|2009ApJ...694..222C|1 sigma|        61 GHz       | Broad-band measurement|00 47 25 -25 16 00 (J2000)| Flux integrated from map|                                        |From new raw data
187|61 GHz (WMAP)       | 1.0       |+/-0.10 |Jy                  |6.10E+10|  1.00E+00|+/-1.00E-01|Jy|2011ApJS..192...15G|uncertainty|        61 GHz       | Broad-band measurement|00 47 20 -25 13 (J2000)| Flux integrated from map|                                        |From new raw data
188|V (WMAP)            | 1.0       |+/-0.20 | Jy                 |6.10E+10|  1.00E+00|+/-2.00E-01|Jy|2009ApJS..180..283W|uncertainty|        61 GHz       | Broad-band measurement|00 47 19 -25 14 00 (J2000)| Flux integrated from map|                                        |From new raw data
189|41 GHz (WMAP)       | 1164      |+/-184  | milliJy            |4.10E+10|  1.16E+00|+/-1.84E-01|Jy|2009MNRAS.392..733M|uncertainty|        41 GHz       | Broad-band measurement|011.9206 -25.2878 (J2000)| Flux integrated from map|                                        |From new raw data
190|41 GHz (WMAP)       | 1100      ||milliJy             |4.10E+10|  1.10E+00||Jy|2009A&A...508..107G|no uncertainty reported|        41 GHz       | Broad-band measurement|00 47 33.1 -25 17 17.0 (J2000)| Flux integrated from map|                                        |From new raw data
191|41 GHz (WMAP)       | 1.0       |+/-0.2  |Jy                  |4.10E+10|  1.00E+00|+/-2.00E-01|Jy|2009ApJ...694..222C|1 sigma|        41 GHz       | Broad-band measurement|00 47 25 -25 16 00 (J2000)| Flux integrated from map|                                        |From new raw data
192|Q (WMAP)            | 1.1       |+/-0.10 | Jy                 |4.10E+10|  1.10E+00|+/-1.00E-01|Jy|2009ApJS..180..283W|uncertainty|        41 GHz       | Broad-band measurement|00 47 19 -25 14 00 (J2000)| Flux integrated from map|                                        |From new raw data
193|41 GHz (WMAP)       | 1.1       |+/-0.09 |Jy                  |4.10E+10|  1.10E+00|+/-9.00E-02|Jy|2011ApJS..192...15G|uncertainty|        41 GHz       | Broad-band measurement|00 47 20 -25 13 (J2000)| Flux integrated from map|                                        |From new raw data
194|41 GHz (WMAP)       | 1.3       |+/-0.3  |Jy                  |4.10E+10|  1.30E+00|+/-3.00E-01|Jy|2003ApJS..148...97B|uncertainty|      41   GHz       | Broad-band measurement|004717.7 -251228 (J2000)| Flux integrated from map|                                        |From new raw data
195|33 GHz (WMAP)       | 985       |+/-193  | milliJy            |3.30E+10|  9.85E-01|+/-1.93E-01|Jy|2009MNRAS.392..733M|uncertainty|        33 GHz       | Broad-band measurement|011.9206 -25.2878 (J2000)| Flux integrated from map|                                        |From new raw data
196|33 GHz (WMAP)       | 0.9       |+/-0.09 |Jy                  |3.30E+10|  9.00E-01|+/-9.00E-02|Jy|2011ApJS..192...15G|uncertainty|        33 GHz       | Broad-band measurement|00 47 20 -25 13 (J2000)| Flux integrated from map|                                        |From new raw data
197|33 GHz (WMAP)       | 0.4       |+/-0.2  |Jy                  |3.30E+10|  4.00E-01|+/-2.00E-01|Jy|2003ApJS..148...97B|uncertainty|      33   GHz       | Broad-band measurement|004717.7 -251228 (J2000)| Flux integrated from map|                                        |From new raw data
198|33 GHz (EVLA)       | 314.27    |+/-0.05 |milliJy             |3.30E+10|  3.14E-01|+/-5.00E-05|Jy|2011ApJ...739L..24K|uncertainty|    33.0   GHz       | Broad-band measurement|| Flux integrated from map|                                        |From new raw data
199|Ka (WMAP)           | 0.9       |+/-0.10 | Jy                 |3.30E+10|  9.00E-01|+/-1.00E-01|Jy|2009ApJS..180..283W|uncertainty|        33 GHz       | Broad-band measurement|00 47 19 -25 14 00 (J2000)| Flux integrated from map|                                        |From new raw data
200|H58{alpha} (EVLA)   | 44.3E-22  |+/-0.7E-22|W/m^2^              |3.29E+10|  4.43E+05|+/-7.00E+03|Jy-Hz|2011ApJ...739L..24K|uncertainty|    32.852 GHz       | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|                                        |From new raw data
201|32 GHz (EVLA)       | 332.5     |+/-0.1  |milliJy             |3.20E+10|  3.33E-01|+/-1.00E-04|Jy|2011ApJ...739L..24K|uncertainty|    32.0   GHz       | Broad-band measurement|| Flux integrated from map|                                        |From new raw data
202|31400 MHz           | 0.59      |+/-.08  |Jy                  |3.14E+10|  5.90E-01|+/-8.00E-02|Jy|1981AJ.....86.1306G|uncertainty|   31400   MHz       | Broad-band measurement|004505.50 -253341.0 (B1950)| Not reported in paper|From Kuhr catalog (1981A&AS...45..367K) |Transformed from previously published data
203|H59{alpha} (EVLA)   | 39.9E-22  |+/-0.8E-22|W/m^2^              |3.12E+10|  3.99E+05|+/-8.00E+03|Jy-Hz|2011ApJ...739L..24K|uncertainty|    31.223 GHz       | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|                                        |From new raw data
204|23 GHz (WMAP)       | 1097      |+/-157  | milliJy            |2.30E+10|  1.10E+00|+/-1.57E-01|Jy|2009MNRAS.392..733M|uncertainty|        23 GHz       | Broad-band measurement|011.9206 -25.2878 (J2000)| Flux integrated from map|                                        |From new raw data
205|23 GHz (WMAP)       | 1.2       |+/-0.05 |Jy                  |2.30E+10|  1.20E+00|+/-5.00E-02|Jy|2011ApJS..192...15G|uncertainty|        23 GHz       | Broad-band measurement|00 47 20 -25 13 (J2000)| Flux integrated from map|                                        |From new raw data
206|23 GHz (WMAP)       | 1.3       |+/-0.1  |Jy                  |2.30E+10|  1.30E+00|+/-1.00E-01|Jy|2003ApJS..148...97B|uncertainty|      23   GHz       | Broad-band measurement|004717.7 -251228 (J2000)| Flux integrated from map|                                        |From new raw data
207|K (WMAP)            | 1.1       |+/-0.06 | Jy                 |2.30E+10|  1.10E+00|+/-6.00E-02|Jy|2009ApJS..180..283W|uncertainty|        23 GHz       | Broad-band measurement|00 47 19 -25 14 00 (J2000)| Flux integrated from map|                                        |From new raw data
208|23 GHz (VLA)        | 0.56      |+/-0.06 |Jy                  |2.30E+10|  5.60E-01|+/-6.00E-02|Jy|2005PASJ...57..549T|uncertainty|      23   GHz       | Broad-band measurement|| Total flux|                                        |From new raw data
209|22 GHz (ATCA)       | 0.489     |+/-0.049|Jy                  |2.20E+10|  4.89E-01|+/-4.90E-02|Jy|2006A&A...445..465R|uncertainty|      22   GHz       | Broad-band measurement|| Modelled datum|                                        |From new raw data
210|20 GHz (ATCA)       | 608       |+/-29   |milliJy             |1.99E+10|  6.08E-01|+/-2.90E-02|Jy|2010MNRAS.402.2403M|rms uncertainty|    19.904 GHz       | Broad-band measurement|00 47 33.08 -25 17 17.7 (J2000)| Flux integrated from map|Flux may be unreliable                  |From new raw data
211|18.5 GHz (ATCA)     | 0.571     |+/-0.029|Jy                  |1.85E+10|  5.71E-01|+/-2.90E-02|Jy|2006A&A...445..465R|uncertainty|    18.5   GHz       | Broad-band measurement|| Modelled datum|                                        |From new raw data
212|10695 MHz           | 0.87      |+/-.06  |Jy                  |1.07E+10|  8.70E-01|+/-6.00E-02|Jy|1981A&AS...45..367K|uncertainty|   10695   MHz       | Broad-band measurement|004505.50 -253341.0 (B1950)| Not reported in paper|                                        |From new raw data
213|8870 MHz            | 1.47      |+/-.06  |Jy                  |8.87E+09|  1.47E+00|+/-6.00E-02|Jy|1973AuJPh..26...93S|uncertainty|    8870   MHz       | Broad-band measurement|004505.50 -253341.0 (B1950)| Not reported in paper|From Kuhr catalog (1981A&AS...45..367K) |Transformed from previously published data
214|8400 MHz            | 1.26      ||Jy                  |8.40E+09|  1.26E+00||Jy|1990PKS90.C...0000W|no uncertainty reported|    8400   MHz       | Broad-band measurement|00 45 05.7 -25 33 40 (B1950)| Integrated from scans|                                        |Homogenized from new and previously published data
215|3.6 cm (Effelsberg) | 980       |+/-50   | milliJy            |8.35E+09|  9.80E-01|+/-5.00E-02|Jy|2009A&A...494..563H|uncertainty|       3.6 cm        | Broad-band measurement|00 47 33.12 -25 17 17.3 (J2000)| Total flux|                                        |From new raw data
216|8 GHz (ATCA)        | 1411      |+/-34   |milliJy             |8.00E+09|  1.41E+00|+/-3.40E-02|Jy|2010MNRAS.402.2403M|rms uncertainty|         8 GHz       | Broad-band measurement|00 47 33.08 -25 17 17.7 (J2000)| Flux integrated from map|Flux may be unreliable                  |From new raw data
217|7.0 GHz (ATA)       | 1.55      |+/-0.09 |Jy                  |7.00E+09|  1.55E+00|+/-9.00E-02|Jy|2010ApJ...710.1462W|uncertainty|       7.0 GHz       | Broad-band measurement|| Flux integrated from map|Total flux; Calibrator is 3C 147        |From new raw data
218|7.0 GHz (ATA)       | 1.04      |+/-0.04 |Jy                  |7.00E+09|  1.04E+00|+/-4.00E-02|Jy|2010ApJ...710.1462W|uncertainty|       7.0 GHz       | Broad-band measurement|| Flux integrated from map|Core flux; Calibrator is 3C 147         |From new raw data
219|6.7 GHz (ATA)       | 1.87      |+/-0.15 |Jy                  |6.70E+09|  1.87E+00|+/-1.50E-01|Jy|2010ApJ...710.1462W|uncertainty|       6.7 GHz       | Broad-band measurement|| Flux integrated from map|Total flux; Calibrator is 3C 147        |From new raw data
220|6.7 GHz (ATA)       | 1.13      |+/-0.04 |Jy                  |6.70E+09|  1.13E+00|+/-4.00E-02|Jy|2010ApJ...710.1462W|uncertainty|       6.7 GHz       | Broad-band measurement|| Flux integrated from map|Core flux; Calibrator is 3C 147         |From new raw data
221|6.4 GHz (ATA)       | 1.18      |+/-0.04 |Jy                  |6.40E+09|  1.18E+00|+/-4.00E-02|Jy|2010ApJ...710.1462W|uncertainty|       6.4 GHz       | Broad-band measurement|| Flux integrated from map|Core flux; Calibrator is 3C 147         |From new raw data
222|6.4 GHz (ATA)       | 1.72      |+/-0.09 |Jy                  |6.40E+09|  1.72E+00|+/-9.00E-02|Jy|2010ApJ...710.1462W|uncertainty|       6.4 GHz       | Broad-band measurement|| Flux integrated from map|Total flux; Calibrator is 3C 147        |From new raw data
223|6.3 GHz (ATA)       | 1.16      |+/-0.03 |Jy                  |6.30E+09|  1.16E+00|+/-3.00E-02|Jy|2010ApJ...710.1462W|uncertainty|       6.3 GHz       | Broad-band measurement|| Flux integrated from map|Core flux; Calibrator is 3C 147         |From new raw data
224|6.3 GHz (ATA)       | 1.68      |+/-0.08 |Jy                  |6.30E+09|  1.68E+00|+/-8.00E-02|Jy|2010ApJ...710.1462W|uncertainty|       6.3 GHz       | Broad-band measurement|| Flux integrated from map|Total flux; Calibrator is 3C 147        |From new raw data
225|6.1 GHz (ATA)       | 1.76      |+/-0.07 |Jy                  |6.10E+09|  1.76E+00|+/-7.00E-02|Jy|2010ApJ...710.1462W|uncertainty|       6.1 GHz       | Broad-band measurement|| Flux integrated from map|Total flux; Calibrator is 3C 147        |From new raw data
226|6.1 GHz (ATA)       | 1.16      |+/-0.03 |Jy                  |6.10E+09|  1.16E+00|+/-3.00E-02|Jy|2010ApJ...710.1462W|uncertainty|       6.1 GHz       | Broad-band measurement|| Flux integrated from map|Core flux; Calibrator is 3C 147         |From new raw data
227|6.0 GHz (ATA)       | 1.95      |+/-0.08 |Jy                  |6.00E+09|  1.95E+00|+/-8.00E-02|Jy|2010ApJ...710.1462W|uncertainty|       6.0 GHz       | Broad-band measurement|| Flux integrated from map|Total flux; Calibrator is 3C 147        |From new raw data
228|6.0 GHz (ATA)       | 1.20      |+/-0.03 |Jy                  |6.00E+09|  1.20E+00|+/-3.00E-02|Jy|2010ApJ...710.1462W|uncertainty|       6.0 GHz       | Broad-band measurement|| Flux integrated from map|Core flux; Calibrator is 3C 147         |From new raw data
229|5.9 GHz (ATA)       | 1.21      |+/-0.04 |Jy                  |5.90E+09|  1.21E+00|+/-4.00E-02|Jy|2010ApJ...710.1462W|uncertainty|       5.9 GHz       | Broad-band measurement|| Flux integrated from map|Core flux; Calibrator is 3C 147         |From new raw data
230|5.9 GHz (ATA)       | 1.97      |+/-0.09 |Jy                  |5.90E+09|  1.97E+00|+/-9.00E-02|Jy|2010ApJ...710.1462W|uncertainty|       5.9 GHz       | Broad-band measurement|| Flux integrated from map|Total flux; Calibrator is 3C 147        |From new raw data
231|5.8 GHz (ATA)       | 1.87      |+/-0.08 |Jy                  |5.80E+09|  1.87E+00|+/-8.00E-02|Jy|2010ApJ...710.1462W|uncertainty|       5.8 GHz       | Broad-band measurement|| Flux integrated from map|Total flux; Calibrator is 3C 147        |From new raw data
232|5.8 GHz (ATA)       | 1.26      |+/-0.04 |Jy                  |5.80E+09|  1.26E+00|+/-4.00E-02|Jy|2010ApJ...710.1462W|uncertainty|       5.8 GHz       | Broad-band measurement|| Flux integrated from map|Core flux; Calibrator is 3C 147         |From new raw data
233|5.7 GHz (ATA)       | 1.26      |+/-0.03 |Jy                  |5.70E+09|  1.26E+00|+/-3.00E-02|Jy|2010ApJ...710.1462W|uncertainty|       5.7 GHz       | Broad-band measurement|| Flux integrated from map|Core flux; Calibrator is 3C 147         |From new raw data
234|5.7 GHz (ATA)       | 2.01      |+/-0.09 |Jy                  |5.70E+09|  2.01E+00|+/-9.00E-02|Jy|2010ApJ...710.1462W|uncertainty|       5.7 GHz       | Broad-band measurement|| Flux integrated from map|Total flux; Calibrator is 3C 147        |From new raw data
235|5.6 GHz (ATA)       | 2.20      |+/-0.10 |Jy                  |5.60E+09|  2.20E+00|+/-1.00E-01|Jy|2010ApJ...710.1462W|uncertainty|       5.6 GHz       | Broad-band measurement|| Flux integrated from map|Total flux; Calibrator is 3C 147        |From new raw data
236|5.6 GHz (ATA)       | 1.30      |+/-0.03 |Jy                  |5.60E+09|  1.30E+00|+/-3.00E-02|Jy|2010ApJ...710.1462W|uncertainty|       5.6 GHz       | Broad-band measurement|| Flux integrated from map|Core flux; Calibrator is 3C 147         |From new raw data
237|5.1 GHz (ATA)       | 2.23      |+/-0.17 |Jy                  |5.10E+09|  2.23E+00|+/-1.70E-01|Jy|2010ApJ...710.1462W|uncertainty|       5.1 GHz       | Broad-band measurement|| Flux integrated from map|Total flux; Calibrator is 3C 48         |From new raw data
238|5.1 GHz (ATA)       | 1.34      |+/-0.07 |Jy                  |5.10E+09|  1.34E+00|+/-7.00E-02|Jy|2010ApJ...710.1462W|uncertainty|       5.1 GHz       | Broad-band measurement|| Flux integrated from map|Core flux; Calibrator is 3C 48          |From new raw data
239|5010 MHz            | 2.08      |+/-0.208|Jy                  |5.01E+09|  2.08E+00|+/-2.08E-01|Jy|1970ApL.....5...29W|estimated error|5010       MHz       | Broad-band measurement|| Flux in fixed aperture|                                        |From new raw data
240|5009 MHz            | 2.52      |+/-.23  |Jy                  |5.01E+09|  2.52E+00|+/-2.30E-01|Jy|1981A&AS...45..367K|uncertainty|    5009   MHz       | Broad-band measurement|004505.50 -253341.0 (B1950)| Not reported in paper|Recal. to Baars scale by factor of 1.03 |Recalibrated data
241|5009 MHz            | 2.14      |+/-.09  |Jy                  |5.01E+09|  2.14E+00|+/-9.00E-02|Jy|1981A&AS...45..367K|uncertainty|    5009   MHz       | Broad-band measurement|004505.50 -253341.0 (B1950)| Not reported in paper|Recal. to Baars scale by factor of 1.03 |Recalibrated data
242|5.0 GHz (ATA)       | 1.45      |+/-0.04 |Jy                  |5.00E+09|  1.45E+00|+/-4.00E-02|Jy|2010ApJ...710.1462W|uncertainty|       5.0 GHz       | Broad-band measurement|| Flux integrated from map|Core flux; Calibrator is 3C 147         |From new raw data
243|5.0 GHz (ATA)       | 1.37      |+/-0.10 |Jy                  |5.00E+09|  1.37E+00|+/-1.00E-01|Jy|2010ApJ...710.1462W|uncertainty|       5.0 GHz       | Broad-band measurement|| Flux integrated from map|Core flux; Calibrator is 3C 48          |From new raw data
244|5.0 GHz (ATA)       | 2.01      |+/-0.18 |Jy                  |5.00E+09|  2.01E+00|+/-1.80E-01|Jy|2010ApJ...710.1462W|uncertainty|       5.0 GHz       | Broad-band measurement|| Flux integrated from map|Total flux; Calibrator is 3C 48         |From new raw data
245|5.0 GHz (ATA)       | 2.26      |+/-0.10 |Jy                  |5.00E+09|  2.26E+00|+/-1.00E-01|Jy|2010ApJ...710.1462W|uncertainty|       5.0 GHz       | Broad-band measurement|| Flux integrated from map|Total flux; Calibrator is 3C 147        |From new raw data
246|5 GHz (ATCA)        | 2190      |+/-56   |milliJy             |5.00E+09|  2.19E+00|+/-5.60E-02|Jy|2010MNRAS.402.2403M|rms uncertainty|         5 GHz       | Broad-band measurement|00 47 33.08 -25 17 17.7 (J2000)| Flux integrated from map|Flux may be unreliable                  |From new raw data
247|5000 MHz            | 2.080     ||Jy                  |5.00E+09|  2.08E+00||Jy|1990PKS90.C...0000W|no uncertainty reported|    5000   MHz       | Broad-band measurement|00 45 05.7 -25 33 40 (B1950)| Integrated from scans|                                        |Homogenized from new and previously published data
248|4.9 GHz (ATA)       | 1.35      |+/-0.04 |Jy                  |4.90E+09|  1.35E+00|+/-4.00E-02|Jy|2010ApJ...710.1462W|uncertainty|       4.9 GHz       | Broad-band measurement|| Flux integrated from map|Core flux; Calibrator is 3C 147         |From new raw data
249|4.9 GHz (ATA)       | 2.35      |+/-0.08 |Jy                  |4.90E+09|  2.35E+00|+/-8.00E-02|Jy|2010ApJ...710.1462W|uncertainty|       4.9 GHz       | Broad-band measurement|| Flux integrated from map|Total flux; Calibrator is 3C 147        |From new raw data
250|6.2 cm (Effelsberg) | 1270      |+/-60   | milliJy            |4.85E+09|  1.27E+00|+/-6.00E-02|Jy|2009A&A...494..563H|uncertainty|       6.2 cm        | Broad-band measurement|00 47 33.12 -25 17 17.3 (J2000)| Total flux|                                        |From new raw data
251|4.85 GHz            | 2433      |+/-99   |milliJy             |4.85E+09|  2.43E+00|+/-9.90E-02|Jy|1994ApJS...90..179G|rms noise|4.85       GHz       | Broad-band measurement|004732.4 -251716 (J2000)| Modelled datum|                                        |From new raw data; Corrected for contaminating sources
252|4.8 GHz (Effelsberg)| 2707      ||milliJy             |4.80E+09|  2.71E+00||Jy|2009ApJ...693.1392S|no uncertainty reported|       4.8 GHz       | Broad-band measurement|| Flux integrated from map|                                        |From reprocessed raw data
253|4.7 GHz (ATA)       | 1.47      |+/-0.03 |Jy                  |4.70E+09|  1.47E+00|+/-3.00E-02|Jy|2010ApJ...710.1462W|uncertainty|       4.7 GHz       | Broad-band measurement|| Flux integrated from map|Core flux; Calibrator is 3C 147         |From new raw data
254|4.7 GHz (ATA)       | 2.47      |+/-0.10 |Jy                  |4.70E+09|  2.47E+00|+/-1.00E-01|Jy|2010ApJ...710.1462W|uncertainty|       4.7 GHz       | Broad-band measurement|| Flux integrated from map|Total flux; Calibrator is 3C 147        |From new raw data
255|4.6 GHz (ATA)       | 1.46      |+/-0.04 |Jy                  |4.60E+09|  1.46E+00|+/-4.00E-02|Jy|2010ApJ...710.1462W|uncertainty|       4.6 GHz       | Broad-band measurement|| Flux integrated from map|Core flux; Calibrator is 3C 147         |From new raw data
256|4.6 GHz (ATA)       | 2.51      |+/-0.08 |Jy                  |4.60E+09|  2.51E+00|+/-8.00E-02|Jy|2010ApJ...710.1462W|uncertainty|       4.6 GHz       | Broad-band measurement|| Flux integrated from map|Total flux; Calibrator is 3C 147        |From new raw data
257|4.5 GHz (ATA)       | 2.47      |+/-0.04 |Jy                  |4.50E+09|  2.47E+00|+/-4.00E-02|Jy|2010ApJ...710.1462W|uncertainty|       4.5 GHz       | Broad-band measurement|| Flux integrated from map|Total flux; Calibrator is 3C 147        |From new raw data
258|4.5 GHz (ATA)       | 1.50      |+/-0.02 |Jy                  |4.50E+09|  1.50E+00|+/-2.00E-02|Jy|2010ApJ...710.1462W|uncertainty|       4.5 GHz       | Broad-band measurement|| Flux integrated from map|Core flux; Calibrator is 3C 147         |From new raw data
259|3.7 GHz (ATA)       | 1.75      |+/-0.08 |Jy                  |3.70E+09|  1.75E+00|+/-8.00E-02|Jy|2010ApJ...710.1462W|uncertainty|       3.7 GHz       | Broad-band measurement|| Flux integrated from map|Core flux; Calibrator is 3C 147         |From new raw data
260|3.7 GHz (ATA)       | 2.90      |+/-0.19 |Jy                  |3.70E+09|  2.90E+00|+/-1.90E-01|Jy|2010ApJ...710.1462W|uncertainty|       3.7 GHz       | Broad-band measurement|| Flux integrated from map|Total flux; Calibrator is 3C 147        |From new raw data
261|3.6 GHz (ATA)       | 1.75      |+/-0.04 |Jy                  |3.60E+09|  1.75E+00|+/-4.00E-02|Jy|2010ApJ...710.1462W|uncertainty|       3.6 GHz       | Broad-band measurement|| Flux integrated from map|Core flux; Calibrator is 3C 147         |From new raw data
262|3.6 GHz (ATA)       | 3.13      |+/-0.08 |Jy                  |3.60E+09|  3.13E+00|+/-8.00E-02|Jy|2010ApJ...710.1462W|uncertainty|       3.6 GHz       | Broad-band measurement|| Flux integrated from map|Total flux; Calibrator is 3C 147        |From new raw data
263|3.3 GHz (ATA)       | 1.76      |+/-0.02 |Jy                  |3.30E+09|  1.76E+00|+/-2.00E-02|Jy|2010ApJ...710.1462W|uncertainty|       3.3 GHz       | Broad-band measurement|| Flux integrated from map|Core flux; Calibrator is 3C 147         |From new raw data
264|3.3 GHz (ATA)       | 3.16      |+/-0.04 |Jy                  |3.30E+09|  3.16E+00|+/-4.00E-02|Jy|2010ApJ...710.1462W|uncertainty|       3.3 GHz       | Broad-band measurement|| Flux integrated from map|Total flux; Calibrator is 3C 147        |From new raw data
265|3.1 GHz (ATA)       | 1.83      |+/-0.02 |Jy                  |3.10E+09|  1.83E+00|+/-2.00E-02|Jy|2010ApJ...710.1462W|uncertainty|       3.1 GHz       | Broad-band measurement|| Flux integrated from map|Core flux; Calibrator is 3C 147         |From new raw data
266|3.1 GHz (ATA)       | 3.34      |+/-0.04 |Jy                  |3.10E+09|  3.34E+00|+/-4.00E-02|Jy|2010ApJ...710.1462W|uncertainty|       3.1 GHz       | Broad-band measurement|| Flux integrated from map|Total flux; Calibrator is 3C 147        |From new raw data
267|3.1 GHz (ATA)       | 1.89      |+/-0.06 |Jy                  |3.10E+09|  1.89E+00|+/-6.00E-02|Jy|2010ApJ...710.1462W|uncertainty|       3.1 GHz       | Broad-band measurement|| Flux integrated from map|Core flux; Calibrator is 3C 48          |From new raw data
268|3.1 GHz (ATA)       | 3.59      |+/-0.11 |Jy                  |3.10E+09|  3.59E+00|+/-1.10E-01|Jy|2010ApJ...710.1462W|uncertainty|       3.1 GHz       | Broad-band measurement|| Flux integrated from map|Total flux; Calibrator is 3C 48         |From new raw data
269|3.0 GHz (ATA)       | 1.98      |+/-0.07 |Jy                  |3.00E+09|  1.98E+00|+/-7.00E-02|Jy|2010ApJ...710.1462W|uncertainty|       3.0 GHz       | Broad-band measurement|| Flux integrated from map|Core flux; Calibrator is 3C 48          |From new raw data
270|3.0 GHz (ATA)       | 3.74      |+/-0.12 |Jy                  |3.00E+09|  3.74E+00|+/-1.20E-01|Jy|2010ApJ...710.1462W|uncertainty|       3.0 GHz       | Broad-band measurement|| Flux integrated from map|Total flux; Calibrator is 3C 48         |From new raw data
271|2700 MHz            | 3.520     ||Jy                  |2.70E+09|  3.52E+00||Jy|1990PKS90.C...0000W|no uncertainty reported|    2700   MHz       | Broad-band measurement|00 45 05.7 -25 33 40 (B1950)| Integrated from scans|                                        |Homogenized from new and previously published data
272|2.7 GHz (ATA)       | 3.75      |+/-0.04 |Jy                  |2.70E+09|  3.75E+00|+/-4.00E-02|Jy|2010ApJ...710.1462W|uncertainty|       2.7 GHz       | Broad-band measurement|| Flux integrated from map|Total flux; Calibrator is 3C 147        |From new raw data
273|2.7 GHz (ATA)       | 2.01      |+/-0.02 |Jy                  |2.70E+09|  2.01E+00|+/-2.00E-02|Jy|2010ApJ...710.1462W|uncertainty|       2.7 GHz       | Broad-band measurement|| Flux integrated from map|Core flux; Calibrator is 3C 147         |From new raw data
274|2700 MHz            | 3.52      |+/-.12  |Jy                  |2.70E+09|  3.52E+00|+/-1.20E-01|Jy|1976AuJPA..39....1W|uncertainty|    2700   MHz       | Broad-band measurement|004505.50 -253341.0 (B1950)| Not reported in paper|From Kuhr catalog (1981A&AS...45..367K) |Transformed from previously published data
275|2695 MHz            | 3.72      |+/-.05  |Jy                  |2.70E+09|  3.72E+00|+/-5.00E-02|Jy|1981A&AS...45..367K|uncertainty|    2695   MHz       | Broad-band measurement|004505.50 -253341.0 (B1950)| Not reported in paper|Recal. to Baars scale by factor of 1.011|Recalibrated data
276|2650 MHz            | 3.88      |+/-.12  |Jy                  |2.65E+09|  3.88E+00|+/-1.20E-01|Jy|1975AuJPA..38....1W|uncertainty|    2650   MHz       | Broad-band measurement|004505.50 -253341.0 (B1950)| Not reported in paper|From Kuhr catalog (1981A&AS...45..367K) |Transformed from previously published data
277|2.6 GHz (ATA)       | 1.95      |+/-0.03 |Jy                  |2.60E+09|  1.95E+00|+/-3.00E-02|Jy|2010ApJ...710.1462W|uncertainty|       2.6 GHz       | Broad-band measurement|| Flux integrated from map|Core flux; Calibrator is 3C 147         |From new raw data
278|2.6 GHz (ATA)       | 3.75      |+/-0.06 |Jy                  |2.60E+09|  3.75E+00|+/-6.00E-02|Jy|2010ApJ...710.1462W|uncertainty|       2.6 GHz       | Broad-band measurement|| Flux integrated from map|Total flux; Calibrator is 3C 147        |From new raw data
279|2.1 GHz (ATA)       | 2.25      |+/-0.08 |Jy                  |2.10E+09|  2.25E+00|+/-8.00E-02|Jy|2010ApJ...710.1462W|uncertainty|       2.1 GHz       | Broad-band measurement|| Flux integrated from map|Core flux; Calibrator is 3C 48          |From new raw data
280|2.1 GHz (ATA)       | 4.21      |+/-0.12 |Jy                  |2.10E+09|  4.21E+00|+/-1.20E-01|Jy|2010ApJ...710.1462W|uncertainty|       2.1 GHz       | Broad-band measurement|| Flux integrated from map|Total flux; Calibrator is 3C 48         |From new raw data
281|2.0 GHz (ATA)       | 4.64      |+/-0.12 |Jy                  |2.00E+09|  4.64E+00|+/-1.20E-01|Jy|2010ApJ...710.1462W|uncertainty|       2.0 GHz       | Broad-band measurement|| Flux integrated from map|Total flux; Calibrator is 3C 48         |From new raw data
282|2.0 GHz (ATA)       | 2.35      |+/-0.08 |Jy                  |2.00E+09|  2.35E+00|+/-8.00E-02|Jy|2010ApJ...710.1462W|uncertainty|       2.0 GHz       | Broad-band measurement|| Flux integrated from map|Core flux; Calibrator is 3C 48          |From new raw data
283|1.9 GHz (ATA)       | 4.78      |+/-0.08 |Jy                  |1.90E+09|  4.78E+00|+/-8.00E-02|Jy|2010ApJ...710.1462W|uncertainty|       1.9 GHz       | Broad-band measurement|| Flux integrated from map|Total flux; Calibrator is 3C 147        |From new raw data
284|1.9 GHz (ATA)       | 2.36      |+/-0.05 |Jy                  |1.90E+09|  2.36E+00|+/-5.00E-02|Jy|2010ApJ...710.1462W|uncertainty|       1.9 GHz       | Broad-band measurement|| Flux integrated from map|Core flux; Calibrator is 3C 147         |From new raw data
285|1.8 GHz (ATA)       | 2.39      |+/-0.05 |Jy                  |1.80E+09|  2.39E+00|+/-5.00E-02|Jy|2010ApJ...710.1462W|uncertainty|       1.8 GHz       | Broad-band measurement|| Flux integrated from map|Core flux; Calibrator is 3C 147         |From new raw data
286|1.8 GHz (ATA)       | 4.89      |+/-0.08 |Jy                  |1.80E+09|  4.89E+00|+/-8.00E-02|Jy|2010ApJ...710.1462W|uncertainty|       1.8 GHz       | Broad-band measurement|| Flux integrated from map|Total flux; Calibrator is 3C 147        |From new raw data
287|1.7 GHz (ATA)       | 2.48      |+/-0.05 |Jy                  |1.70E+09|  2.48E+00|+/-5.00E-02|Jy|2010ApJ...710.1462W|uncertainty|       1.7 GHz       | Broad-band measurement|| Flux integrated from map|Core flux; Calibrator is 3C 147         |From new raw data
288|1.7 GHz (ATA)       | 5.16      |+/-0.09 |Jy                  |1.70E+09|  5.16E+00|+/-9.00E-02|Jy|2010ApJ...710.1462W|uncertainty|       1.7 GHz       | Broad-band measurement|| Flux integrated from map|Total flux; Calibrator is 3C 147        |From new raw data
289|1.5 GHz (ATA)       | 5.13      |+/-0.13 |Jy                  |1.50E+09|  5.13E+00|+/-1.30E-01|Jy|2010ApJ...710.1462W|uncertainty|       1.5 GHz       | Broad-band measurement|| Flux integrated from map|Total flux; Calibrator is 3C 48         |From new raw data
290|1.5 GHz (ATA)       | 2.54      |+/-0.08 |Jy                  |1.50E+09|  2.54E+00|+/-8.00E-02|Jy|2010ApJ...710.1462W|uncertainty|       1.5 GHz       | Broad-band measurement|| Flux integrated from map|Core flux; Calibrator is 3C 48          |From new raw data
291|HI (21 cm line)     | 9.57      |+/-0.10 |m_21 mag            |1.42E+09|  6.49E+06|+/-6.26E+05|Jy-Hz|1991RC3.9.C...0000d|rms uncertainty|21         cm        | Line measurement; flux integrated over line; lines measured in emission|004505.7 -253340 (B1950)| Multiple methods|m_21 equiv. to S(HI) = 6.486E-20 W m^-2 |Homogenized from new and previously published data
292|HI 21 cm line       | 834.85    ||Jy km s^-1^         |1.42E+09|  3.95E+06||Jy-Hz|2005ApJS..160..149S|no uncertainty reported|242        km s^-1^  | Line measurement; flux integrated over line; lines measured in emission|00 47 34.9 -25 17 17 (J2000)| Flux integrated from map|Corrected line flux                     |From new raw data
293|HI line (Parkes)    | 693.5     ||Jy km s^-1^         |1.42E+09|  3.28E+06||Jy-Hz|2005MNRAS.361...34D|no uncertainty reported|258.8      km s^-1^  | Line measurement; flux integrated over line; lines measured in emission|004731.1 -251723. (J2000)| Flux integrated from map|                                        |Averaged from previously published data
294|HI 21 cm line       | 544.54    ||Jy km s^-1^         |1.42E+09|  2.58E+06||Jy-Hz|2005ApJS..160..149S|no uncertainty reported|242        km s^-1^  | Line measurement; flux integrated over line; lines measured in emission|00 47 34.9 -25 17 17 (J2000)| Flux integrated from map|                                        |From new raw data
295|HI 21cm line Parkes | 692.9     |+/-42.2 | Jy km/s            |1.42E+09|  3.27E+06|+/-1.99E+05|Jy-Hz|2004AJ....128...16K|uncertainty|     243   km s^-1^  | Line measurement; flux integrated over line|00 47 31 -25 17 22 (J2000)| Flux integrated from map|Extended source                         |From new raw data
296|HI 21 cm line       | 999.99    |+/-152.24|Jy km s^-1^         |1.42E+09|  4.73E+06|+/-7.20E+05|Jy-Hz|2005ApJS..160..149S|uncertainty|242        km s^-1^  | Line measurement; flux integrated over line; lines measured in emission|00 47 34.9 -25 17 17 (J2000)| Flux integrated from map|Self-absorption corrected line flux     |From new raw data
297|HI (21 cm line)     | 924.80    ||Jy km s^-1^         |1.42E+09|  4.36E+06||Jy-Hz|1989H&RHI.C...0000H|no uncertainty reported|21         cm        | Line measurement; flux integrated over line; lines measured in emission|004507.6 -253339. (B1950)| Not reported in paper|                                        |Transformed from previously published data
298|HI (21 cm line)     ||<380.00    |Jy km s^-1^         |1.42E+09||1.80E+06|Jy-Hz|1989H&RHI.C...0000H|no uncertainty reported|21         cm        | Line measurement; flux integrated over line; not detected|004507.6 -253339. (B1950)| Not reported in paper|                                        |Transformed from previously published data
299|HI (21 cm line)     | 756.30    |+/-74.30|Jy km s^-1^         |1.42E+09|  3.57E+06|+/-3.50E+05|Jy-Hz|1989H&RHI.C...0000H|no uncertainty reported|21         cm        | Line measurement; flux integrated over line; lines measured in emission|004507.6 -253339. (B1950)| Not reported in paper|                                        |Transformed from previously published data
300|HI (21 cm line)     | 1429.00   ||Jy km s^-1^         |1.42E+09|  6.74E+06||Jy-Hz|1989H&RHI.C...0000H|no uncertainty reported|21         cm        | Line measurement; flux integrated over line; lines measured in emission|004507.6 -253339. (B1950)| Not reported in paper|                                        |Transformed from previously published data
301|HI (21 cm line)     | 794.60    |+/-8.90 |Jy km s^-1^         |1.42E+09|  3.75E+06|+/-4.20E+04|Jy-Hz|1989H&RHI.C...0000H|no uncertainty reported|21         cm        | Line measurement; flux integrated over line; lines measured in emission|004507.6 -253339. (B1950)| Not reported in paper|                                        |Transformed from previously published data
302|1410 MHz            | 6.18      |+/-.12  |Jy                  |1.41E+09|  6.18E+00|+/-1.20E-01|Jy|1981A&AS...45..367K|uncertainty|    1410   MHz       | Broad-band measurement|004505.50 -253341.0 (B1950)| Not reported in paper|Recal. to Baars scale by factor of 1.017|Recalibrated data
303|1410 MHz            | 6.000     ||Jy                  |1.41E+09|  6.00E+00||Jy|1990PKS90.C...0000W|no uncertainty reported|    1410   MHz       | Broad-band measurement|00 45 05.7 -25 33 40 (B1950)| Integrated from scans|                                        |Homogenized from new and previously published data
304|1.4GHz              | 2994.7    |+/-113.5|milliJy             |1.40E+09|  3.00E+00|+/-1.14E-01|Jy|1998AJ....115.1693C|uncertainty|    1.40   GHz       | Broad-band measurement|00 47 33.13 -25 17 17.1 (J2000)| Flux integrated from map|High Integral                           |From new raw data
305|1.4 GHz (ATA)       | 2.76      |+/-0.09 |Jy                  |1.40E+09|  2.76E+00|+/-9.00E-02|Jy|2010ApJ...710.1462W|uncertainty|       1.4 GHz       | Broad-band measurement|| Flux integrated from map|Core flux; Calibrator is 3C 48          |From new raw data
306|1.4 GHz (ATA)       | 5.97      |+/-0.09 |Jy                  |1.40E+09|  5.97E+00|+/-9.00E-02|Jy|2010ApJ...710.1462W|uncertainty|       1.4 GHz       | Broad-band measurement|| Flux integrated from map|Total flux; Calibrator is 3C 147        |From new raw data
307|1.4 GHz (ATA)       | 5.93      |+/-0.13 |Jy                  |1.40E+09|  5.93E+00|+/-1.30E-01|Jy|2010ApJ...710.1462W|uncertainty|       1.4 GHz       | Broad-band measurement|| Flux integrated from map|Total flux; Calibrator is 3C 48         |From new raw data
308|1.4 GHz (ATA)       | 2.75      |+/-0.06 |Jy                  |1.40E+09|  2.75E+00|+/-6.00E-02|Jy|2010ApJ...710.1462W|uncertainty|       1.4 GHz       | Broad-band measurement|| Flux integrated from map|Core flux; Calibrator is 3C 147         |From new raw data
309|1.4 GHz (VLA)       | 5704.5    || milliJy            |1.40E+09|  5.70E+00||Jy|2004ApJ...606..829S|no uncertainty reported|     1.4   GHz       | Broad-band measurement|00 47 33.2 -25 17 16.2 (J2000)| Total flux|                                        |From reprocessed raw data
310|1.3 GHz (ATA)       | 6.29      |+/-0.07 |Jy                  |1.30E+09|  6.29E+00|+/-7.00E-02|Jy|2010ApJ...710.1462W|uncertainty|       1.3 GHz       | Broad-band measurement|| Flux integrated from map|Total flux; Calibrator is 3C 147        |From new raw data
311|1.3 GHz (ATA)       | 2.78      |+/-0.04 |Jy                  |1.30E+09|  2.78E+00|+/-4.00E-02|Jy|2010ApJ...710.1462W|uncertainty|       1.3 GHz       | Broad-band measurement|| Flux integrated from map|Core flux; Calibrator is 3C 147         |From new raw data
312|1.2 GHz (ATA)       | 6.75      |+/-0.10 |Jy                  |1.20E+09|  6.75E+00|+/-1.00E-01|Jy|2010ApJ...710.1462W|uncertainty|       1.2 GHz       | Broad-band measurement|| Flux integrated from map|Total flux; Calibrator is 3C 147        |From new raw data
313|1.2 GHz (ATA)       | 2.93      |+/-0.05 |Jy                  |1.20E+09|  2.93E+00|+/-5.00E-02|Jy|2010ApJ...710.1462W|uncertainty|       1.2 GHz       | Broad-band measurement|| Flux integrated from map|Core flux; Calibrator is 3C 147         |From new raw data
314|1.1 GHz (ATA)       | 2.98      |+/-0.05 |Jy                  |1.10E+09|  2.98E+00|+/-5.00E-02|Jy|2010ApJ...710.1462W|uncertainty|       1.1 GHz       | Broad-band measurement|| Flux integrated from map|Core flux; Calibrator is 3C 147         |From new raw data
315|1.1 GHz (ATA)       | 6.90      |+/-0.08 |Jy                  |1.10E+09|  6.90E+00|+/-8.00E-02|Jy|2010ApJ...710.1462W|uncertainty|       1.1 GHz       | Broad-band measurement|| Flux integrated from map|Total flux; Calibrator is 3C 147        |From new raw data
316|960 MHz             | 8.1       |+/-.12  |Jy                  |9.60E+08|  8.10E+00|+/-1.20E-01|Jy|1981A&AS...45..367K|uncertainty|     960   MHz       | Broad-band measurement|004505.50 -253341.0 (B1950)| Not reported in paper|Recal. to Baars scale by factor of 1.029|Recalibrated data
317|635 MHz             | 10.87     |+/-.25  |Jy                  |6.35E+08|  1.09E+01|+/-2.50E-01|Jy|1981A&AS...45..367K|uncertainty|     635   MHz       | Broad-band measurement|004505.50 -253341.0 (B1950)| Not reported in paper|Recal. to Baars scale by factor of 1.035|Recalibrated data
318|468 MHz             | 15.17     |+/-1.54 |Jy                  |4.68E+08|  1.52E+01|+/-1.54E+00|Jy|1981A&AS...45..367K|uncertainty|     468   MHz       | Broad-band measurement|004505.50 -253341.0 (B1950)| Not reported in paper|Recal. to Baars scale by factor of 1.045|Recalibrated data
319|408 MHz             | 6.120     ||Jy                  |4.08E+08|  6.12E+00||Jy|1990PKS90.C...0000W|no uncertainty reported|     408   MHz       | Broad-band measurement|00 45 05.7 -25 33 40 (B1950)| Integrated from scans|                                        |Homogenized from new and previously published data
320|408 MHz             | 6.12      |+/-0.29 |Jy                  |4.08E+08|  6.12E+00|+/-2.90E-01|Jy|1981MNRAS.194..693L|rms noise|408        MHz       | Broad-band measurement|004505.6 -253337 (B1950)| Modelled datum|Extended source; flux density may be low|From new raw data; Corrected for contaminating sources
321|365 MHz (Texas)     | 3.350     |+/-0.139|Jy                  |3.65E+08|  3.35E+00|+/-1.39E-01|Jy|1996AJ....111.1945D|internal error|365        MHz       | Broad-band measurement; obtained by interpolation over frequency|004505.750 -253339.80 (B1950)| Integrated from scans|Model:D;MFlag:+;EFlag:+;LFlag:+.        |From new raw data
322|160 MHz             | 11.9      ||Jy                  |1.60E+08|  1.19E+01||Jy|1995AuJPh..48..143S|no uncertainty reported|160        MHz       | Broad-band measurement|004505.2 -253353. (B1950)| Flux integrated from map|                                        |From new raw data
323|145 MHz (PAPER)     | 13.1      ||Jy                  |1.45E+08|  1.31E+01||Jy|2011ApJ...734L..34J|no uncertainty reported|       145 MHz       | Broad-band measurement|11.95 -25.37 (J2000)| Flux integrated from map|                                        |From new raw data
324|80 MHz              | 25.       ||Jy                  |8.00E+07|  2.50E+01||Jy|1995AuJPh..48..143S|no uncertainty reported| 80        MHz       | Broad-band measurement|004505.2 -253353. (B1950)| Flux integrated from map|                                        |From new raw data
325|80 MHz              | 24        |+/-4.00 |Jy                  |8.00E+07|  2.40E+01|+/-4.00E+00|Jy|1981A&AS...45..367K|uncertainty|      80   MHz       | Broad-band measurement|004505.50 -253341.0 (B1950)| Not reported in paper|Recal. to Baars scale by factor of 1.074|Recalibrated data
326|80 MHz              | 22.00     ||Jy                  |8.00E+07|  2.20E+01||Jy|1990PKS90.C...0000W|no uncertainty reported|      80   MHz       | Broad-band measurement|00 45 05.7 -25 33 40 (B1950)| Integrated from scans|                                        |Homogenized from new and previously published data
327|74 MHz (VLA)        | 10.87     |+/-1.12 | Jy                 |7.38E+07|  1.09E+01|+/-1.12E+00|Jy|2007AJ....134.1245C|rms uncertainty|    73.8   MHz       | Broad-band measurement|00 47 33.42 -25 17 13.9 (J2000)| Flux integrated from map|Corrected for clean bias                |From new raw data
328|57.5 MHz            | 48.0      |+/-9.0  |Jy                  |5.75E+07|  4.80E+01|+/-9.00E+00|Jy|1990ApJ...352...30I|uncertainty|57.5       MHz       | Broad-band measurement|| Flux integrated from map|                                        |From new raw data
