
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-04-05T08:15:36PDT



Photometric Data for SDSS J163655.77+405910.0

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|24 microns (MIPS)   | 473.0     |57      |mJy             |1.27E+13|473.E-03|+/-57.E-03|Jy|2009ApJ...694.1517D|3sigma uncertainty|     23.68 microns   | Broad-band measurement|12 37 11.89 +62 22 11.8 (J2000)| Flux integrated from map|                                        |From new raw data
2|70 microns (MIPS)   | 1.4       |+/-0.4  |mJy             |4.20E+12|1.4E-03|0.4E-03|Jy|2009ApJ...699.1610H|3 sigma|     71.42 microns   | Broad-band measurement|221804.42 +002154.4 (J2000)| Flux in fixed aperture|                                        |From new raw data
3|350 microns (SHARC-II) |           |<36.0   |mJy             |8.565E+11|      |36.0E-03|Jy|2005MNRAS.358..149P|3sigma uncertainty|     850   microns   | Broad-band measurement|12 37 11.7 +62 22 12 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
4|850 microns (SCUBA) |           |<3.6    |mJy             |3.53E+11|  |3.6E-03|Jy|2005MNRAS.358..149P|3rms uncertainty|     850   microns   | Broad-band measurement|12 37 11.7 +62 22 12 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
5|1200 microns (MAMBO)|           |<6.6    |mJy             |2.50E+11|  |6.6E-03|Jy|2004MNRAS.354..779G|3rms uncertainty|      1200 microns   | Broad-band measurement|16 36 55.9 +40 59 12 (J2000)| Flux integrated from map|S/N = 3.66                              |From new raw data
6|1.4 GHz (VLA)       | 126.3     |+/-8.6  | microJy        |1.40E+09| 126.3E-06|+/-8.6E-06|Jy|2006MNRAS.371..963B|1 sigma|       1.4 GHz       | Broad-band measurement|16 36 55.767 +40 59 09.97 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
