
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-06-14T16:33:23PDT



Photometric Data for [HB89] 1623+269:MD0066

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|G (WHT)             | 24.32     ||mag                 |6.38E+14|  6.79E-07||Jy|2006ApJ...647..128E|no uncertainty reported|    0.47   microns   | Broad-band measurement|| Flux in fixed aperture|                                        |Averaged from previously published data
5|J (Hale/WIRC)       | 21.89     ||mag                 |2.40E+14|  2.74E-06||Jy|2006ApJ...646..107E|no uncertainty reported|    1.25   microns   | Broad-band measurement|16 25 40.39 +26 50 08.88 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data; derived from aflux in a different band and a color
6|K_s (Hale/WIRC)     | 20.15     ||mag                 |1.39E+14|  5.84E-06||Jy|2006ApJ...646..107E|no uncertainty reported|    2.15   microns   | Broad-band measurement|16 25 40.39 +26 50 08.88 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data
