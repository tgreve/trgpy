
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-04-05T08:15:36PDT



Photometric Data for SDSS J163655.77+405910.0

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|R (Subaru)          | 24.0      |+/-0.3  |mag                 |4.76E+14|  7.84E-07|+/-2.17E-07|Jy|2006ApJS..167..103F|rms uncertainty|    6300   A         | Broad-band measurement|| Flux in fixed aperture|3" radius aperture                      |From new raw data
2|I (Cousins)         | 24.15     |+/-0.14 |mag                 |3.79E+14|  5.58E-07|+/-7.68E-08|Jy|2004ApJ...616...71S|1 sigma|    7900   A         | Broad-band measurement|| Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
3|z (Subaru)          | 23.1      |+/-0.5  |mag                 |3.26E+14|  1.26E-06|+/-5.80E-07|Jy|2006ApJS..167..103F|rms uncertainty|    9200   A         | Broad-band measurement|| Flux in fixed aperture|3" radius aperture                      |From new raw data
4|J (2MASS)           | 21.53     |+/-0.19 |mag                 |2.40E+14|  3.89E-06|+/-7.44E-07|Jy|2004ApJ...616...71S|1 sigma|    1.25   microns   | Broad-band measurement|| Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
5|K_s (2MASS)         | 19.36     |+/-0.10 |mag                 |1.38E+14|  1.20E-05|+/-1.16E-06|Jy|2004ApJ...616...71S|1 sigma|    2.17   microns   | Broad-band measurement|| Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
1|24 microns (MIPS)   | 105.0     |15      |microJy             |1.27E+13|105.E-06|+/-15.E-06|Jy|2009ApJ...694.1517D|3sigma uncertainty|     23.68 microns   | Broad-band measurement|12 37 11.89 +62 22 11.8 (J2000)| Flux integrated from map|                                        |From new raw data
2|850 microns (SCUBA) |           |<5.7    |mJy             |3.53E+11|  |5.7E-03|Jy|2005MNRAS.358..149P|3sigma uncertainty|     850   microns   | Broad-band measurement|12 37 11.7 +62 22 12 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
3|1.4 GHz (VLA)       |     44.9  |+/-2.4  |uJy             |1.40E+09| 44.9E-06|+/-2.4E-06|Jy|2006MNRAS.371..963B|1 sigma|       1.4 GHz       | Broad-band measurement|16 36 55.767 +40 59 09.97 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
7|1.4 GHz (VLA)       | 61        |+/-10   |microJy             |1.40E+09|  6.10E-05|+/-1.00E-05|Jy|2006ApJS..167..103F|uncertainty|     1.4   GHz       | Broad-band measurement|13 12 07.737 +42 39 44.92 (J2000)| Flux integrated from map|Corrected to the sky; see paper         |From new raw data
