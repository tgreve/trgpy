
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-05-28T01:50:15PDT



Photometric Data for PJ020941.3, z=2.5534

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
4|UKIDSS J            | 0.04   |+/-0.001|mJy        |2.40161e+14|0.04E-3|+/-0.001E-3|Jy|2010Natur.464..733S|3rms uncertainty reported|      3344 A         | Broad-band measurement|21 35 11.6 -01 02 52.0 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
5|UKIDSS H            | 0.06   |+/-0.01|mJy         |1.83775e+14|0.06E-3|+/-0.01E-3|Jy|2010Natur.464..733S|3rms uncertainty reported|      3344 A         | Broad-band measurement|21 35 11.6 -01 02 52.0 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
6|UKIDSS K            | 0.05   |+/-0.01|mJy         |1.36207e+14|0.05E-3|+/-0.01E-3|Jy|2010Natur.464..733S|3rms uncertainty reported|      3344 A         | Broad-band measurement|21 35 11.6 -01 02 52.0 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
1|3.4 microns (WISE)  | 1.22      |+/-0.03|mJy          |8.82E+13|  1.22E-03|+/-0.03E-03|Jy|2012AJ....144...49W|uncertainty|       3.4 microns   | Broad-band measurement|213.942657 +11.495400 (J2000)| Not reported in paper|                                        |Averaged from previously published data
2|4.6 microns (WISE)  | 1.30      |+/-0.03|mJy          |6.52E+13|  1.30E-03|+/-0.03E-03|Jy|2012AJ....144...49W|uncertainty|       4.6 microns   | Broad-band measurement|213.942657 +11.495400 (J2000)| Not reported in paper|                                        |Averaged from previously published data
3|12 microns (WISE)   | 0.61      |+/-0.12|mJy          |2.50E+13|  0.61E-03|+/-0.12E-03|Jy|2012AJ....144...49W|uncertainty|        12 microns   | Broad-band measurement|213.942657 +11.495400 (J2000)| Not reported in paper|                                        |Averaged from previously published data
4|22 microns (WISE)   | 4.35      |+/-0.87|mJy          |1.36E+13|  4.35E-03|+/-0.87E-03|Jy|2012AJ....144...49W|uncertainty|        22 microns   | Broad-band measurement|213.942657 +11.495400 (J2000)| Not reported in paper|                                        |Averaged from previously published data
1|250 microns (SPIRE) | 824.0     |+/-82.  |mJy         |1.199e+12|824.0E-03 |+/-82.0e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
1|250 microns (SPIRE) | 826.0     |+/-7.  |mJy         |1.199e+12|826.0E-03 |+/-7.0e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
3|350 microns (SPIRE) | 897.0     |+/-89.  |mJy         |8.565e+11|897.0E-03 |+/-89.0e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
3|350 microns (SPIRE) | 912.0     |+/-7.  |mJy         |8.565e+11|912.0E-03 |+/-7.0e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
5|350 microns (PLANCK) | 877.0    |+/-375.  |mJy        |8.55e+11|877.0E-03 |+/-375.0e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
17|450 microns (SCUBA) | 217.0    |+/-72. |milliJy      |6.66E+11|  217.E-03|+/-72.E-03 |Jy|2002MNRAS.331..495S|no uncertainty reported|     450   microns   | Broad-band measurement|140105.0 +025225 (J2000)| Flux integrated from map|                                        |From new raw data
5|500 microns (SPIRE) | 703.0     |+/-70.  |mJy         |5.996e+11|703.0E-03 |+/-70.0e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
5|500 microns (SPIRE) | 717.0     |+/-8.  |mJy         |5.996e+11|717.0E-03 |+/-8.0e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
9|850 microns (SCUBA) | 167.0     |+/-4. |milliJy       |3.53E+11|  167.E-03|+/-4.E-03 |Jy|2002MNRAS.331..495S|no uncertainty reported|     850   microns   | Broad-band measurement|140105.0 +025225 (J2000)| Flux integrated from map|                                        |From new raw data
2|1.1mm (AzTEC)        | 147. |+/-15.| mJy  | 2.73E11| 147.E-3| 15.E-3 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
2|1.1mm (AzTEC)        | 95.5 |+/-2.4| mJy  | 2.73E11| 95.5E-3| 2.4E-3 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
5|VLA Ka-band 33.8GHz  |  244   |+/-38 |mJy          |33.8372E+9|244.0E-06 |+/-38E-06|Jy|2010ApJ...709..210K|uncertainty|      870  microns   | Broad-band measurement|16 35 55.67 +66 12 59.51 (J2000)| Flux integrated from map|                                        |From new raw data
5|VLA K-band 22.0GHz    |  200   |+/-51 |mJy          |21.999E+9|200.0E-06 |+/-51E-06|Jy|2010ApJ...709..210K|uncertainty|      870  microns   | Broad-band measurement|16 35 55.67 +66 12 59.51 (J2000)| Flux integrated from map|                                        |From new raw data
14|5.0GHz (VLA)        | 1000.0    |+/- 300. |uJy  | 5.0E9   | 1000.E-6|+/-300.E-6 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
14|1.4GHz (VLA)        | 1595.    |+/-342 |uJy  | 1.4E9   | 1595.E-6|+/-342.E-6 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
14|1.4GHz (VLA)        | 3.23    |+/-0.121 |uJy  | 1.4E9   | 3.23E-3|+/-0.121E-3 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
14|1.4GHz (VLA)        | 2.15    |+/-0.121 |uJy  | 1.4E9   | 2.15E-3|+/-0.121E-3 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
