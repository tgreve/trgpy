
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-04-04T05:13:41PDT



Photometric Data for Bolocam LE 1100.08

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|B (SUBARU) AB       | 26.45     |+/-0.09 | mag                |6.69E+14|  9.55E-08|+/-7.92E-09|Jy|2008MNRAS.386.1107D|uncertainty|      4478 A         | Broad-band measurement|10 52 38.299 +57 24 35.76 (J2000)| Flux in fixed aperture|3" diameter aperture                    |From new raw data
2|R (SUBARU)          | 24.34     |+/-0.05 |mag                 |4.68E+14|  5.66E-07|+/-2.60E-08|Jy|2005MNRAS.364.1025I|uncertainty|    6400   A         | Broad-band measurement| | Flux in fixed aperture|                                        |Averaged new and previously published data
3|R (SUBARU) AB       | 24.90     |+/-0.06 | mag                |4.58E+14|  3.98E-07|+/-2.20E-08|Jy|2008MNRAS.386.1107D|uncertainty|      6550 A         | Broad-band measurement|10 52 38.299 +57 24 35.76 (J2000)| Flux in fixed aperture|3" diameter aperture                    |From new raw data
4|I (Cousins)         | 23.26     |+/-0.16 |mag                 |3.79E+14|  1.27E-06|+/-2.01E-07|Jy|2004ApJ...616...71S|1 sigma|    7900   A         | Broad-band measurement| | Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
5|I (SUBARU) AB       | 24.21     |+/-0.06 | mag                |3.75E+14|  7.52E-07|+/-4.15E-08|Jy|2008MNRAS.386.1107D|uncertainty|      7996 A         | Broad-band measurement|10 52 38.299 +57 24 35.76 (J2000)| Flux in fixed aperture|3" diameter aperture                    |From new raw data
6|z (SUBARU) AB       | 23.47     |+/-0.06 | mag                |3.31E+14|  1.49E-06|+/-8.21E-08|Jy|2008MNRAS.386.1107D|uncertainty|      9054 A         | Broad-band measurement|10 52 38.299 +57 24 35.76 (J2000)| Flux in fixed aperture|3" diameter aperture                    |From new raw data
7|F160W (HST) AB      | 22.43     |+/-0.08 |mag                 |1.87E+14|  3.87E-06|+/-2.85E-07|Jy|2010MNRAS.405..234S|uncertainty|      1.60 microns   | Broad-band measurement|10 52 38.30 +57 24 35.8 (J2000)| Flux in fixed aperture|                                        |From new raw data
8|K_s_ (2MASS)        | 20.32     |+/-0.24 |mag                 |1.38E+14|  4.97E-06|+/-1.23E-06|Jy|2004ApJ...616...71S|1 sigma|    2.17   microns   | Broad-band measurement| | Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
9|K (UKIRT) AB        | 21.39     |+/-0.06 | mag                |1.36E+14|  1.01E-05|+/-5.58E-07|Jy|2008MNRAS.386.1107D|uncertainty|      2.20 microns   | Broad-band measurement|10 52 38.299 +57 24 35.76 (J2000)| Flux in fixed aperture|3" diameter aperture                    |From new raw data
10|3.6 microns IRAC AB | 20.66     |+/-0.21 | mag                |8.44E+13|  1.98E-05|+/-3.82E-06|Jy|2008MNRAS.386.1107D|uncertainty|     3.550 microns   | Broad-band measurement|10 52 38.299 +57 24 35.76 (J2000)| Flux in fixed aperture|3" diameter aperture                    |From new raw data
11|3.6 microns (IRAC)  | 29.7      |+/-3.2  |microJy             |8.44E+13|  2.97E-05|+/-3.20E-06|Jy|2009ApJ...699.1610H|uncertainty|     3.550 microns   | Broad-band measurement|10 52 38.30 +57 24 35.7 (J2000)| Flux in fixed aperture|                                        |From new raw data
12|4.5 microns IRAC AB | 20.67     |+/-0.20 | mag                |6.67E+13|  1.96E-05|+/-3.61E-06|Jy|2008MNRAS.386.1107D|uncertainty|     4.493 microns   | Broad-band measurement|10 52 38.299 +57 24 35.76 (J2000)| Flux in fixed aperture|3" diameter aperture                    |From new raw data
13|4.5 microns (IRAC)  | 33.6      |+/-3.6  |microJy             |6.67E+13|  3.36E-05|+/-3.60E-06|Jy|2009ApJ...699.1610H|uncertainty|     4.493 microns   | Broad-band measurement|10 52 38.30 +57 24 35.7 (J2000)| Flux in fixed aperture|                                        |From new raw data
14|5.8 microns IRAC AB | 20.47     |+/-0.39 | mag                |5.23E+13|  2.36E-05|+/-8.46E-06|Jy|2008MNRAS.386.1107D|uncertainty|     5.731 microns   | Broad-band measurement|10 52 38.299 +57 24 35.76 (J2000)| Flux in fixed aperture|3" diameter aperture                    |From new raw data
15|5.8 microns (IRAC)  | 30.7      |+/-4.7  |microJy             |5.23E+13|  3.07E-05|+/-4.70E-06|Jy|2009ApJ...699.1610H|uncertainty|     5.731 microns   | Broad-band measurement|10 52 38.30 +57 24 35.7 (J2000)| Flux in fixed aperture|                                        |From new raw data
18|8.0 microns (IRAC)  | |<58.8      |microJy             |3.85E+13| |5.88E-05|Jy|2009ApJ...699.1610H|3 sigma|     7.782 microns   | Broad-band measurement|10 52 38.30 +57 24 35.7 (J2000)| Flux in fixed aperture|                                        |From new raw data
19|8.0 microns IRAC AB | 21.09     |+/-0.44 | mag                |3.81E+13|  1.33E-05|+/-5.39E-06|Jy|2008MNRAS.386.1107D|uncertainty|     7.872 microns   | Broad-band measurement|10 52 38.299 +57 24 35.76 (J2000)| Flux in fixed aperture|3" diameter aperture                    |From new raw data
20|PAH 8.6 (Spitzer)   | 0.52E-15  |+/-0.16E-15|erg/s/cm^2^         |3.49E+13|  1.49E-06|+/-4.58E-07|Jy|2009ApJ...699..667M|rms uncertainty|       8.6 microns   | Line measurement; flux integrated over line; lines measured in emission|10 52 38.30 +57 24 35.8 (J2000)| Flux integrated from map|                                        |From new raw data
21|24 microns (Spitzer)| 175.0     |+/-23.0 | microJy            |1.27E+13|  1.75E-04|+/-2.30E-05|Jy|2007MNRAS.380..199I|rms uncertainty|     23.68 microns   | Broad-band measurement|10 52 38.31 +57 24 34.8 (J2000)| Flux integrated from map|                                        |Averaged from previously published data
22|24 microns (MIPS)   | 322.0     |+/-38.0 |microJy             |1.27E+13|  3.22E-04|+/-3.80E-05|Jy|2009ApJ...699.1610H|uncertainty|     23.68 microns   | Broad-band measurement|105238.30 +572435.8 (J2000)| Flux in fixed aperture|                                        |From new raw data
23|70 microns (MIPS)   | |<6.4       |milliJy             |4.20E+12| |6.40E-03|Jy|2009ApJ...699.1610H|3 sigma|     71.42 microns   | Broad-band measurement|105238.30 +572435.8 (J2000)| Flux in fixed aperture|                                        |From new raw data
24|350 microns (CSO)   | 40.5      |+/-6.5  | milliJy            |8.57E+11|  4.05E-02|+/-6.50E-03|Jy|2008MNRAS.384.1597C|uncertainty|       350 microns   | Broad-band measurement| | Flux integrated from map|Corrected for flux boosting             |From new raw data
25|350 microns (SHARC2)| 40.5      |+/-6.5  |milliJy             |8.57E+11|  4.05E-02|+/-6.50E-03|Jy|2006ApJ...650..592K|uncertainty|     350   microns   | Broad-band measurement| | Total flux|                                        |From new raw data
26|850 microns (SCUBA) | 10.9      |+/-2.4  |milliJy             |3.53E+11|  1.09E-02|+/-2.40E-03|Jy|2005ApJ...622..772C|uncertainty|     850   microns   | Broad-band measurement|105238.30 +572435.8 (J2000)| Flux integrated from map|                                        |From new raw data
27|850 microns (SCUBA) | 11.0      |+/-2.3  |mag                 |3.53E+11|  1.10E-02|+/-2.30E-03|Jy|2006MNRAS.370.1057S|uncertainty|     850   microns   | Broad-band measurement|10 52 38.21 +57 24 35.1 (J2000)| From fitting to map|S/N = 5.33                              |From reprocessed raw data
28|850 microns (SCUBA) | 10.9      |+/-1.9  | milliJy            |3.53E+11|  1.09E-02|+/-1.90E-03|Jy|2007MNRAS.380..199I|rms uncertainty|       850 microns   | Broad-band measurement|10 52 38.247 +57 24 36.54 (J2000)| Flux integrated from map|                                        |Averaged from previously published data
29|0.85 mm (SCUBA)     | 10.9      |+/-2.1  |milliJy             |3.53E+11|  1.09E-02|+/-2.10E-03|Jy|2005MNRAS.364.1025I|uncertainty|    0.85   mm        | Broad-band measurement|105238.6 +572438 (J2000)| Flux integrated from map|                                        |Averaged from previously published data
31|1.2 mm (MAMBO)      | 4.8       |+/-0.6  |milliJy             |2.50E+11|  4.80E-03|+/-6.00E-04|Jy|2005MNRAS.364.1025I|uncertainty|     1.2   mm        | Broad-band measurement|105238.3 +572437 (J2000)| Flux integrated from map|                                        |Averaged from previously published data
32|1200 microns (MAMBO)| 4.8       |+/-0.6  | milliJy            |2.50E+11|  4.80E-03|+/-6.00E-04|Jy|2004MNRAS.354..779G|uncertainty|      1200 microns   | Broad-band measurement|10 52 38.3 +57 24 37 (J2000)| Flux integrated from map|S/N = 8.00                              |From new raw data
33|1.4 GHz (VLA)       | 35.0      |+/-5.2  | microJy            |1.40E+09|  3.50E-05|+/-5.20E-06|Jy|2007MNRAS.380..199I|rms uncertainty|       1.4 GHz       | Broad-band measurement|10 52 38.401 +57 24 39.50 (J2000)| Flux integrated from map|                                        |From reprocessed raw data
34|1.4 GHz (VLA)       | 25.8      |+/-4.9  | microJy            |1.40E+09|  2.58E-05|+/-4.90E-06|Jy|2007MNRAS.380..199I|rms uncertainty|       1.4 GHz       | Broad-band measurement|10 52 38.299 +57 24 35.76 (J2000)| Flux integrated from map|                                        |From reprocessed raw data
35|1.4 GHz (VLA)       | 29        |+/-11   |microJy             |1.40E+09|  2.90E-05|+/-1.10E-05|Jy|2005MNRAS.364.1025I|uncertainty|     1.4   GHz       | Broad-band measurement|105238.30 +572435.8 (J2000)| Flux integrated from map|                                        |Averaged from previously published data
