
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2017-01-03T07:44:13PST



Photometric Data for B2 0748+27

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|CO (8-7) line (IRAM)| 2.2       |+/-0.7  | Jy km/s            |9.24E+11|  1.61E+06|+/-5.14E+05|Jy-Hz|2007A&A...470...53A|uncertainty|    3.1999           | Line measurement; flux integrated over line|| From fitting to map|                                        |From new raw data
2|350 microns (CSO)   | 36        |+/-16   |milliJy             |8.57E+11|  3.60E-02|+/-1.60E-02|Jy|2009ApJ...707..988W|rms noise|       350 microns   | Broad-band measurement|07 51 47.46 +27 16 31.4 (J2000)| Flux integrated from map|S/N=2.3 sigma                           |From new raw data
3|CO (4-3) line (IRAM)| 4.2       |+/-0.7  | Jy km/s            |4.62E+11|  1.54E+06|+/-2.57E+05|Jy-Hz|2007A&A...470...53A|uncertainty|    3.1999           | Line measurement; flux integrated over line|| From fitting to map|                                        |From new raw data
4|CO (3-2) line (IRAM)| 4.6       |+/-0.5  | Jy km/s            |3.44E+11|  1.26E+06|+/-1.37E+05|Jy-Hz|2007A&A...470...53A|uncertainty|    3.1999           | Line measurement; flux integrated over line|| From fitting to map|                                        |From new raw data
5|220 GHz (IRAM/PdBI) | 4.3       |+/-0.8  | milliJy            |2.20E+11|  4.30E-03|+/-8.00E-04|Jy|2007A&A...470...53A|uncertainty|       220 GHz       | Broad-band measurement|| From fitting to map|                                        |From new raw data
6|H_2O (3_13-2_20) VLA||<0.18      |milliJy             |1.83E+11||1.80E-04|Jy|2006ApJ...649..635R|no uncertainty reported|183.3101   GHz       | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|                                        |From new raw data
7|CO(1-0) (EVLA)      | 0.494     |+/-0.105|Jy km/s             |1.15E+11|  4.53E+04|+/-9.61E+03|Jy-Hz|2011ApJ...739L..32R|uncertainty|   115.271 GHz       | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|                                        |From new raw data
8|CO(1-0) (GBT)       | 0.550     |+/-0.095|Jy km/s             |1.15E+11|  5.04E+04|+/-8.70E+03|Jy-Hz|2011ApJ...739L..32R|uncertainty|   115.271 GHz       | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|Measured with Spectrometer backend      |From new raw data
9|110 GHz (IRAM/PdBI) | 3.0       |+/-0.5  | milliJy            |1.10E+11|  3.00E-03|+/-5.00E-04|Jy|2007A&A...470...53A|uncertainty|       110 GHz       | Broad-band measurement|| From fitting to map|                                        |From new raw data
10|82 GHz (IRAM/PdBI)  | 5.1       |+/-0.4  | milliJy            |8.20E+10|  5.10E-03|+/-4.00E-04|Jy|2007A&A...470...53A|uncertainty|        82 GHz       | Broad-band measurement|| From fitting to map|                                        |From new raw data
11|8085 MHz            | 0.12      |+/-0.01 |Jy                  |8.08E+09|  1.20E-01|+/-1.25E-02|Jy|1983AJ.....88...20C|rms uncertainty|8085       MHz       | Broad-band measurement|074837.21 +272415.0 (B1950)| Flux integrated from map|                                        |From new raw data
12|4.85 GHz            | 214       |+/-28   |milliJy             |4.85E+09|  2.14E-01|+/-2.80E-02|Jy|1991ApJS...75.1011G|rms noise|4.85       GHz       | Broad-band measurement|074837.8 +272434 (B1950)| Modelled datum|                                        |From new raw data; Corrected for contaminating sources
13|4.85 GHz            | 209       |+/-15  %|milliJy             |4.85E+09|  2.09E-01|+/-3.14E-02|Jy|1991ApJS...75....1B|uncertainty|4.85       GHz       | Broad-band measurement|074837.9 +272434 (B1950)| Peak flux|                                        |From new raw data; Corrected for contaminating sources
14|4830 MHz (NRAO/GBT)     | 202       ||milliJy             |4.83E+09|  2.02E-01||Jy|1990ApJS...72..621L|no uncertainty reported|    4830   MHz       | Broad-band measurement|07 51 42.0 +27 16 39 (J2000)| Flux integrated from map|S/N = 28                                |From new raw data
15|2695 MHz            | 0.32      |+/-0.02 |Jy                  |2.70E+09|  3.20E-01|+/-1.51E-02|Jy|1983AJ.....88...20C|rms uncertainty|2695       MHz       | Broad-band measurement|074837.21 +272415.0 (B1950)| Flux integrated from map|                                        |From new raw data
16|1.40 GHz (VLA)      | 554       ||milliJy             |1.40E+09|  5.54E-01||Jy|1992ApJS...79..331W|no uncertainty reported|1.4        GHz       | Broad-band measurement|074837.9 +272434 (B1950)| Peak flux|                                        |From new raw data
17|1400 MHz (VLA)      | 0.75      |+/-0.04 |Jy                  |1.40E+09|  7.50E-01|+/-3.81E-02|Jy|1983AJ.....88...20C|rms uncertainty|1400       MHz       | Broad-band measurement|074837.21 +272415.0 (B1950)| Flux integrated from map|                                        |From reprocessed raw data
18|1.4GHz (VLA)        | 595.3     |+/-17.9 |milliJy             |1.40E+09|  5.95E-01|+/-1.79E-02|Jy|1998AJ....115.1693C|uncertainty|    1.40   GHz       | Broad-band measurement|07 51 41.49 +27 16 31.8 (J2000)| Flux integrated from map|                                        |From new raw data
19|408 MHz             | 1.261     |+/-8   %|Jy                  |4.08E+08|  1.26E+00|+/-1.01E-01|Jy|1972A&AS....7....1C|internal error|408        MHz       | Broad-band measurement; peak value reported|074836.9 +272424. (B1950)| Peak flux|                                        |From new raw data
20|365 MHz (Texas)     | 1.469     |+/-0.075|Jy                  |3.65E+08|  1.47E+00|+/-7.50E-02|Jy|1996AJ....111.1945D|internal error|365        MHz       | Broad-band measurement; obtained by interpolation over frequency|074837.099 272416.07 (B1950)| Integrated from scans|Model:D;MFlag:+;EFlag:+;LFlag:+.        |From new raw data
21|74 MHz (VLA)        | 0.89      |+/-0.12 | Jy                 |7.38E+07|  8.90E-01|+/-1.20E-01|Jy|2007AJ....134.1245C|rms uncertainty|    73.8   MHz       | Broad-band measurement|07 51 41.48 +27 16 31.0 (J2000)| Flux integrated from map|Corrected for clean bias                |From new raw data
