
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-04-04T04:53:44PDT



Photometric Data for Bolocam LE 1100.05

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|B (SUBARU) AB       | 24.32     |+/-0.06 | mag                |6.69E+14|  6.79E-07|+/-3.75E-08|Jy|2008MNRAS.386.1107D|uncertainty|      4478 A         | Broad-band measurement|10 52 30.717 +57 22 09.56 (J2000)| Flux in fixed aperture|3" diameter aperture                    |From new raw data
2|R (SUBARU)          | 22.78     |+/-0.02 |mag                 |4.68E+14|  2.38E-06|+/-4.38E-08|Jy|2005MNRAS.364.1025I|uncertainty|    6400   A         | Broad-band measurement| | Flux in fixed aperture|                                        |Averaged new and previously published data
3|R (SUBARU) AB       | 23.74     |+/-0.06 | mag                |4.58E+14|  1.16E-06|+/-6.40E-08|Jy|2008MNRAS.386.1107D|uncertainty|      6550 A         | Broad-band measurement|10 52 30.717 +57 22 09.56 (J2000)| Flux in fixed aperture|3" diameter aperture                    |From new raw data
4|H{alpha} (Keck)     | 1.2E-19   |+/-0.3E-19| W/m^2^             |4.57E+14|  2.63E-08|+/-6.56E-09|Jy|2004ApJ...617...64S|uncertainty|      6563 A         | Line measurement; flux integrated over line; lines measured in emission|105230.73 +572209.5 (J2000)| Flux integrated from map|                                        |From new raw data
5|H{alpha} (IRTF)     | 1.2E-19   |+/-0.5E-19| W/m^2^             |4.57E+14|  2.63E-08|+/-1.09E-08|Jy|2004ApJ...617...64S|uncertainty|      6563 A         | Line measurement; flux integrated over line; lines measured in emission|105230.73 +572209.5 (J2000)| Flux integrated from map|                                        |From new raw data
6|I (Cousins)         | 22.71     |+/-0.07 |mag                 |3.79E+14|  2.10E-06|+/-1.40E-07|Jy|2004ApJ...616...71S|1 sigma|    7900   A         | Broad-band measurement| | Flux in fixed aperture|4" aper; phot contam by near neighbor   |Averaged new and previously published data
7|I (SUBARU) AB       | 23.40     |+/-0.06 | mag                |3.75E+14|  1.59E-06|+/-8.76E-08|Jy|2008MNRAS.386.1107D|uncertainty|      7996 A         | Broad-band measurement|10 52 30.717 +57 22 09.56 (J2000)| Flux in fixed aperture|3" diameter aperture                    |From new raw data
8|z (SUBARU) AB       | 23.18     |+/-0.06 | mag                |3.31E+14|  1.94E-06|+/-1.07E-07|Jy|2008MNRAS.386.1107D|uncertainty|      9054 A         | Broad-band measurement|10 52 30.717 +57 22 09.56 (J2000)| Flux in fixed aperture|3" diameter aperture                    |From new raw data
9|F160W (HST) AB      | 22.11     |+/-0.05 |mag                 |1.87E+14|  5.20E-06|+/-2.39E-07|Jy|2010MNRAS.405..234S|uncertainty|      1.60 microns   | Broad-band measurement|10 52 30.73 +57 22 09.5 (J2000)| Flux in fixed aperture|                                        |From new raw data
10|K_s_ (2MASS)        | 19.22     |+/-0.16 |mag                 |1.38E+14|  1.37E-05|+/-2.17E-06|Jy|2004ApJ...616...71S|1 sigma|    2.17   microns   | Broad-band measurement| | Flux in fixed aperture|4" aper; phot contam by near neighbor   |Averaged new and previously published data
11|K (UKIRT) AB        | 21.06     |+/-0.06 | mag                |1.36E+14|  1.37E-05|+/-7.56E-07|Jy|2008MNRAS.386.1107D|uncertainty|      2.20 microns   | Broad-band measurement|10 52 30.717 +57 22 09.56 (J2000)| Flux in fixed aperture|3" diameter aperture                    |From new raw data
12|3.6 microns IRAC AB | 20.20     |+/-0.19 | mag                |8.44E+13|  3.02E-05|+/-5.29E-06|Jy|2008MNRAS.386.1107D|uncertainty|     3.550 microns   | Broad-band measurement|10 52 30.717 +57 22 09.56 (J2000)| Flux in fixed aperture|3" diameter aperture                    |From new raw data
13|3.6 microns (IRAC)  | 34.3      |+/-3.7  |microJy             |8.44E+13|  3.43E-05|+/-3.70E-06|Jy|2009ApJ...699.1610H|uncertainty|     3.550 microns   | Broad-band measurement|10 52 30.72 +57 22 09.4 (J2000)| Flux in fixed aperture|                                        |From new raw data
14|4.5 microns IRAC AB | 20.15     |+/-0.21 | mag                |6.67E+13|  3.16E-05|+/-6.12E-06|Jy|2008MNRAS.386.1107D|uncertainty|     4.493 microns   | Broad-band measurement|10 52 30.717 +57 22 09.56 (J2000)| Flux in fixed aperture|3" diameter aperture                    |From new raw data
15|4.5 microns (IRAC)  | 40.6      |+/-4.1  |microJy             |6.67E+13|  4.06E-05|+/-4.10E-06|Jy|2009ApJ...699.1610H|uncertainty|     4.493 microns   | Broad-band measurement|10 52 30.72 +57 22 09.4 (J2000)| Flux in fixed aperture|                                        |From new raw data
16|5.8 microns IRAC AB | 20.15     |+/-0.66 | mag                |5.23E+13|  3.16E-05|+/-1.92E-05|Jy|2008MNRAS.386.1107D|uncertainty|     5.731 microns   | Broad-band measurement|10 52 30.717 +57 22 09.56 (J2000)| Flux in fixed aperture|3" diameter aperture                    |From new raw data
17|5.8 microns (IRAC)  | 58.0      |+/-6.7  |microJy             |5.23E+13|  5.80E-05|+/-6.70E-06|Jy|2009ApJ...699.1610H|uncertainty|     5.731 microns   | Broad-band measurement|10 52 30.72 +57 22 09.4 (J2000)| Flux in fixed aperture|                                        |From new raw data
18|8.0 microns (IRAC)  | 47.9      |+/-4.8  |microJy             |3.85E+13|  4.79E-05|+/-4.80E-06|Jy|2009ApJ...699.1610H|uncertainty|     7.782 microns   | Broad-band measurement|10 52 30.72 +57 22 09.4 (J2000)| Flux in fixed aperture|                                        |From new raw data
19|8.0 microns IRAC AB | 20.56     |+/-0.69 | mag                |3.81E+13|  2.17E-05|+/-1.38E-05|Jy|2008MNRAS.386.1107D|uncertainty|     7.872 microns   | Broad-band measurement|10 52 30.717 +57 22 09.56 (J2000)| Flux in fixed aperture|3" diameter aperture                    |From new raw data
20|24 microns (Spitzer)| 188.0     |+/-16.0 | microJy            |1.27E+13|  1.88E-04|+/-1.60E-05|Jy|2007MNRAS.380..199I|rms uncertainty|     23.68 microns   | Broad-band measurement|10 52 30.72 +57 22 09.4 (J2000)| Flux integrated from map|                                        |Averaged from previously published data
21|24 microns (MIPS)   | 177.0     |+/-23.0 |microJy             |1.27E+13|  1.77E-04|+/-2.30E-05|Jy|2009ApJ...699.1610H|uncertainty|     23.68 microns   | Broad-band measurement|105230.73 +572209.5 (J2000)| Flux in fixed aperture|                                        |From new raw data
22|70 microns (MIPS)   | |<4.1       |milliJy             |4.20E+12| |4.10E-03|Jy|2009ApJ...699.1610H|3 sigma|     71.42 microns   | Broad-band measurement|105230.73 +572209.5 (J2000)| Flux in fixed aperture|                                        |From new raw data
23|350 microns (SHARC2)| 41.0      |+/-6.8  |milliJy             |8.57E+11|  4.10E-02|+/-6.80E-03|Jy|2006ApJ...650..592K|uncertainty|     350   microns   | Broad-band measurement| | Total flux|                                        |From new raw data
24|850 microns (SCUBA) | 11        |+/-2.6  |milliJy             |3.53E+11|  1.10E-02|+/-2.60E-03|Jy|2005ApJ...622..772C|uncertainty|     850   microns   | Broad-band measurement|105230.73 +572209.5 (J2000)| Flux integrated from map|                                        |From new raw data
25|0.85 mm (SCUBA)     | 10.8      |+/-2.4  |milliJy             |3.53E+11|  1.08E-02|+/-2.40E-03|Jy|2005MNRAS.364.1025I|uncertainty|    0.85   mm        | Broad-band measurement|105230.4 +572213 (J2000)| Flux integrated from map|                                        |Averaged from previously published data
26|850 microns (SCUBA) | 7.2       |+/-1.9  | milliJy            |3.53E+11|  7.20E-03|+/-1.90E-03|Jy|2007MNRAS.380..199I|rms uncertainty|       850 microns   | Broad-band measurement|10 52 30.110 +57 22 15.55 (J2000)| Flux integrated from map|                                        |Averaged from previously published data
27|850 microns (SCUBA) | 10.8      |+/-2.6  |mag                 |3.53E+11|  1.08E-02|+/-2.60E-03|Jy|2006MNRAS.370.1057S|uncertainty|     850   microns   | Broad-band measurement|10 52 30.39 +57 22 13.2 (J2000)| From fitting to map|S/N = 4.58                              |From reprocessed raw data
28|CO(3-2) line (IRAM) | |<0.6       |Jy km s^-1^         |3.46E+11| |1.55E-07|Jy|2005MNRAS.359.1165G|3 sigma|  2.5901             | Line measurement; flux integrated over line; lines measured in emission|... ... (J2000)| Flux integrated from map|                                        |From new raw data
29|1100 microns (JCMT) | 3.4       |+/-1.0  |milliJy             |2.73E+11|  3.40E-03|+/-1.00E-03|Jy|2010MNRAS.401..160A|uncertainty|      1100 microns   | Broad-band measurement|163.12721 +57.36944 (J2000)| Flux integrated from map|                                        |From new raw data
30|1100 microns (JCMT) | 1.8       |+/-1.0  |milliJy             |2.73E+11|  1.80E-03|+/-1.00E-03|Jy|2010MNRAS.401..160A|uncertainty|      1100 microns   | Broad-band measurement|163.12721 +57.36944 (J2000)| Flux integrated from map|Corrected for boosting                  |From new raw data
31|1.2 mm (MAMBO)      | 2.9       |+/-0.7  |milliJy             |2.50E+11|  2.90E-03|+/-7.00E-04|Jy|2005MNRAS.364.1025I|uncertainty|     1.2   mm        | Broad-band measurement|105229.9 +572205 (J2000)| Flux integrated from map|                                        |Averaged from previously published data
32|1200 microns (MAMBO)| 2.9       |+/-0.7  | milliJy            |2.50E+11|  2.90E-03|+/-7.00E-04|Jy|2004MNRAS.354..779G|uncertainty|      1200 microns   | Broad-band measurement|10 52 29.9 +57 22 05 (J2000)| Flux integrated from map|S/N = 4.14                              |From new raw data
33|1.4 GHz (VLA)       | 54        |+/-14   |microJy             |1.40E+09|  5.40E-05|+/-1.40E-05|Jy|2005MNRAS.364.1025I|uncertainty|     1.4   GHz       | Broad-band measurement|105230.73 +572209.5 (J2000)| Flux integrated from map|                                        |Averaged from previously published data
34|1.4 GHz (VLA)       | 37.4      |+/-4.2  | microJy            |1.40E+09|  3.74E-05|+/-4.20E-06|Jy|2007MNRAS.380..199I|rms uncertainty|       1.4 GHz       | Broad-band measurement|10 52 30.717 +57 22 09.56 (J2000)| Flux integrated from map|                                        |From reprocessed raw data
35|1.4 GHz (VLA)       | 50        |+/-11   | microJy            |1.40E+09|  5.00E-05|+/-1.10E-05|Jy|2006MNRAS.371..963B|1 sigma|       1.4 GHz       | Broad-band measurement|10 52 30.709 +57 22 09.55 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
36|1.4 GHz (VLA)       | 25.3      |+/-4.2  | microJy            |1.40E+09|  2.53E-05|+/-4.20E-06|Jy|2007MNRAS.380..199I|rms uncertainty|       1.4 GHz       | Broad-band measurement|10 52 28.995 +57 22 22.42 (J2000)| Flux integrated from map|                                        |From reprocessed raw data
