
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-06-17T09:40:16PDT



Photometric Data for SDF J132415.7+273058

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
2|i' (Subaru) AB      | 27.56     ||mag                 |3.89E+14|  3.44E-08||Jy|2005PASJ...57..165T|no uncertainty reported|    7709   A         | Broad-band measurement|132408.3 +271543 (J2000)| Flux in fixed aperture|2.0" diam aperture                      |From new raw data
3|z' (Subaru) AB      | 25.96     ||mag                 |3.31E+14|  1.50E-07||Jy|2005PASJ...57..165T|no uncertainty reported|    9054   A         | Broad-band measurement|132408.3 +271543 (J2000)| Flux in fixed aperture|2.0" diam aperture                      |From new raw data
4|NB921 (Subaru) AB   | 24.49     ||mag                 |3.26E+14|  5.81E-07||Jy|2005PASJ...57..165T|no uncertainty reported|    9196   A         | Broad-band measurement|132408.3 +271543 (J2000)| Flux in fixed aperture|2.0" diam aperture                      |From new raw data
5|9500 A (Subaru) AB  | 24.94     ||mag                 |3.16E+14|  3.84E-07||Jy|2005PASJ...57..165T|no uncertainty reported|    9500   A         | Broad-band measurement|132408.3 +271543 (J2000)| Flux in fixed aperture|2.0" diam aperture                      |From new raw data; Corrected for flux in reference beam
11|CARMA 251GHz      |      |<0.75 |mJy                 |2.52E+11|  |0.75E-03|Jy|2011ApJ...736L..28C|1sigma uncertainty|     13006 A         | Broad-band measurement|| Flux in fixed aperture|                                        |From new raw data
