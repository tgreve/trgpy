
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-07-08T08:49:53PDT



Photometric Data for IRAS F08279+5255

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|2-10 keV (ASCA)     | 4.8E-13   ||ergs s^-1^ cm^-2^   |1.45E+18|  3.31E-08||Jy|2005ApJS..161..185U|no uncertainty reported|       6   keV       | Broad-band measurement|127.9283 52.7540 (J2000)| From fitting to map|                                        |From new raw data; Extinction-corrected for Milky Way; NEDfrequency assigned to mid-point of band in keV
2|2-10 keV (Suzaku)   | 4.0E-13   |+/-0.3E-13|erg/cm^2^/s         |1.45E+18|  2.76E-08|+/-2.07E-11|Jy|2009ApJ...697..194S|uncertainty|      6.00 keV       | Broad-band measurement|| Modelled datum|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
3|2-10 keV (XMM)      | 5.0E-13   |+/-0.1E-13|erg/s/cm^2^         |1.45E+18|  3.45E-08|+/-6.90E-10|Jy|2009ApJ...706..644C|uncertainty|      6.00 keV       | Broad-band measurement|| Modelled datum|Absorbed flux                           |From new raw data; NED frequency assigned to mid-point ofband in keV
4|2-10 keV (Chandra)  | 4.5E-13   |+/-0.2E-13|erg/s/cm^2^         |1.45E+18|  3.10E-08|+/-1.38E-09|Jy|2009ApJ...706..644C|uncertainty|      6.00 keV       | Broad-band measurement|| Modelled datum|Absorbed flux                           |From new raw data; NED frequency assigned to mid-point ofband in keV
5|0.3-10 keV (XMM)    | 0.7E-12   ||erg cm^-2^ s^-1^    |1.25E+18|  5.60E-08||Jy|2005MNRAS.364..195P|no uncertainty reported|    5.15   keV       | Broad-band measurement|08 31 41.6 +52 45 17.0 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
6|0.2-10 keV (Chandra)| 6.9E-13   |+/-0.3E-13|erg/cm^2^/s         |1.23E+18|  5.61E-08|+/-2.44E-09|Jy|2008A&A...489...57R|uncertainty|      5.10 keV       | Broad-band measurement|| Modelled datum|                                        |From reprocessed raw data; NED frequency assigned tomid-point of band in keV
7|0.2-10 keV (XMM)    | 7.6E-13   |+/-0.3E-13|erg/cm^2^/s         |1.23E+18|  6.18E-08|+/-2.44E-09|Jy|2008A&A...489...57R|uncertainty|      5.10 keV       | Broad-band measurement|| Modelled datum|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
8|0.5-8 keV (Suzaku)  | 5.63E-13  |+/-0.39E-13|erg/cm^2^/s         |1.03E+18|  5.47E-08|+/-3.79E-09|Jy|2011ApJ...737...91S|uncertainty|      4.25 keV       | Broad-band measurement|| Modelled datum|Obs. date : 2007 Mar 24                 |From reprocessed raw data; Extinction-corrected for MilkyWay; NED frequency assigned to mid-point of band in keV
9|0.5-8 keV (XMM)     | 8.06E-13  |+/-0.15E-13|erg/cm^2^/s         |1.03E+18|  7.83E-08|+/-1.46E-09|Jy|2011ApJ...737...91S|uncertainty|      4.25 keV       | Broad-band measurement|| Modelled datum|Obs. date : 2007 Oct 22                 |From reprocessed raw data; Extinction-corrected for MilkyWay; NED frequency assigned to mid-point of band in keV
10|0.5-8 keV (Chandra) | 5.89E-13  |+/-0.21E-13|erg/cm^2^/s         |1.03E+18|  5.72E-08|+/-2.04E-09|Jy|2011ApJ...737...91S|uncertainty|      4.25 keV       | Broad-band measurement|| Modelled datum|Obs. date : 2008 Jan 14                 |From reprocessed raw data; Extinction-corrected for MilkyWay; NED frequency assigned to mid-point of band in keV
11|0.4-8 keV (Chandra) | 4.7E-13   ||ergs/cm^2^/s        |1.02E+18|  4.61E-08||Jy|2004ApJ...605...45D|no uncertainty reported|    4.20   keV       | Broad-band measurement|| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
12|0.4-8 keV (XMM)     | 5.0E-13   ||ergs/cm^2^/s        |1.02E+18|  4.90E-08||Jy|2004ApJ...605...45D|no uncertainty reported|    4.20   keV       | Broad-band measurement|| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
13|0.7-7 keV (ASCA)    | 5.5E-13   ||ergs s^-1^ cm^-2^   |9.31E+17|  5.91E-08||Jy|2005ApJS..161..185U|no uncertainty reported|    3.85   keV       | Broad-band measurement|127.9283 52.7540 (J2000)| From fitting to map|                                        |From new raw data; Extinction-corrected for Milky Way; NEDfrequency assigned to mid-point of band in keV
14|0.7-2 keV (ASCA)    | 2.0E-13   ||ergs s^-1^ cm^-2^   |3.26E+17|  6.13E-08||Jy|2005ApJS..161..185U|no uncertainty reported|    1.35   keV       | Broad-band measurement|127.9283 52.7540 (J2000)| From fitting to map|                                        |From new raw data; Extinction-corrected for Milky Way; NEDfrequency assigned to mid-point of band in keV
15|0.5-2 keV (Chandra) | 142.9E-15 |+/-2.3E-15| ergs/cm^2^/s       |3.02E+17|  4.73E-08|+/-7.62E-10|Jy|2007ApJ...665.1004J|uncertainty|    1.25   keV       | Broad-band measurement|--- --- (J2000)| Flux integrated from map|                                        |From reprocessed raw data; Extinction-corrected for MilkyWay; NED frequency assigned to mid-point of band in keV
16|0.2-2 keV (XMM)     | 3.5E-13   |+/-0.1E-13|erg/s/cm^2^         |2.66E+17|  1.32E-07|+/-3.76E-09|Jy|2009ApJ...706..644C|uncertainty|      1.10 keV       | Broad-band measurement|| Modelled datum|Absorbed flux                           |From new raw data; NED frequency assigned to mid-point ofband in keV
17|0.2-2 keV (Chandra) | 1.9E-13   |+/-0.2E-13|erg/s/cm^2^         |2.66E+17|  7.14E-08|+/-7.52E-09|Jy|2009ApJ...706..644C|uncertainty|      1.10 keV       | Broad-band measurement|| Modelled datum|Absorbed flux                           |From new raw data; NED frequency assigned to mid-point ofband in keV
18|U (CTIO) AB         | 26.56     || mag                |8.44E+14|  8.63E-08||Jy|2004ApJ...609..513B|no uncertainty reported|      3552 A         | Broad-band measurement|08 31 41.6 +52 45 17 (J2000)| Flux in fixed aperture|3sigma limit                            |From new raw data
19|B (CTIO) AB         | 26.42     || mag                |6.84E+14|  9.82E-08||Jy|2004ApJ...609..513B|no uncertainty reported|      4381 A         | Broad-band measurement|08 31 41.6 +52 45 17 (J2000)| Flux in fixed aperture|3sigma limit                            |From new raw data
20|B (Johnson)         | 18.827    |+/-0.017| mag                |6.81E+14|  1.26E-04|+/-1.97E-06|Jy|2009AJ....138..845O|rms uncertainty|      4400 A         | Broad-band measurement|| Flux in fixed aperture|                                        |From new raw data
21|V (CTIO) AB         | 26.19     || mag                |5.57E+14|  1.21E-07||Jy|2004ApJ...609..513B|no uncertainty reported|   5386.76 A         | Broad-band measurement|08 31 41.6 +52 45 17 (J2000)| Flux in fixed aperture|3sigma limit                            |From new raw data
22|F555W (HST/WFPC2)         | 18.70     |+/-0.07 | mag                |5.54E+14|  1.24E-04|+/-7.96E-06|Jy|2008A&A...478...95Y|uncertainty|      5407 A         | Broad-band measurement|| Modelled datum|                                        |Averaged from previously published data
23|V (Johnson)         | 16.448    |+/-0.012| mag                |5.42E+14|  9.59E-04|+/-1.06E-05|Jy|2009AJ....138..845O|rms uncertainty|      5530 A         | Broad-band measurement|| Flux in fixed aperture|                                        |From new raw data
24|R (JKT)             | 14.5      |+/-0.05 |mag                 |4.58E+14|  4.88E-03|+/-2.25E-04|Jy|2004MNRAS.348..857H|estimated error|    6550   A         | Broad-band measurement|08 31 41.68 +52 45 17.1 (J2000)| Not reported in paper|                                        |From new raw data
25|R (Johnson)         | 15.353    |+/-0.014| mag                |4.33E+14|  2.09E-03|+/-2.69E-05|Jy|2009AJ....138..845O|rms uncertainty|      6930 A         | Broad-band measurement|| Flux in fixed aperture|                                        |From new raw data
26|F814W (HST/WFPC2)         | 16.93     |+/-0.05 | mag                |3.78E+14|  4.21E-04|+/-1.94E-05|Jy|2008A&A...478...95Y|uncertainty|      7940 A         | Broad-band measurement|| Modelled datum|                                        |Averaged from previously published data
27|I (HST)             | 14.55     ||mag                 |3.68E+14|  3.65E-03||Jy|2011ApJ...738...96M|no uncertainty reported|     0.814 microns   | Broad-band measurement|| Not reported in paper|                                        |From reprocessed raw data
28|I (CTIO) AB         | 25.66     || mag                |3.65E+14|  1.98E-07||Jy|2004ApJ...609..513B|no uncertainty reported|   8204.53 A         | Broad-band measurement|08 31 41.6 +52 45 17 (J2000)| Flux in fixed aperture|3sigma limit                            |From new raw data
29|I (JKT)             | 13.9      |+/-0.05 |mag                 |3.63E+14|  7.02E-03|+/-3.23E-04|Jy|2004MNRAS.348..857H|estimated error|    8260   A         | Broad-band measurement|08 31 41.68 +52 45 17.1 (J2000)| Not reported in paper|                                        |From new raw data
30|I (Johnson)         | 14.608    |+/-0.012| mag                |3.41E+14|  3.27E-03|+/-3.62E-05|Jy|2009AJ....138..845O|rms uncertainty|      8785 A         | Broad-band measurement|| Flux in fixed aperture|                                        |From new raw data
31|F160W (HST/NICMOS)         | 15.11     |+/-0.04 | mag                |1.87E+14|  9.43E-04|+/-3.47E-05|Jy|2008A&A...478...95Y|uncertainty|     1.603 microns   | Broad-band measurement|| Modelled datum|                                        |Averaged from previously published data
37|12 microns (IRAS)   ||<1.010E-01 |Jy                  |2.50E+13||1.01E-01|Jy|1990IRASF.C...0000M|90% confidence| 12        microns   | Broad-band measurement|082757.9 +525527 (B1950)| Flux in fixed aperture|                                        |From new raw data
38|3.3 microns Spitzer ||<1.0E-21   | W/cm^2^            |1.85E+13||1.00E+09|Jy-Hz|2004ApJS..154..151S|3 sigma|    16.203 microns   | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|                                        |From new raw data
40|25 microns (IRAS)   | 2.261E-01 |+/-16  %|Jy                  |1.20E+13|  2.26E-01|+/-1.62E-02|Jy|1990IRASF.C...0000M|uncertainty| 25        microns   | Broad-band measurement|082757.9 +525527 (B1950)| Flux in fixed aperture|IRAS quality flag = 2                   |From new raw data
41|6.2 microns Spitzer ||<2.3E-21   | W/cm^2^            |9.85E+12||2.30E+09|Jy-Hz|2004ApJS..154..151S|3 sigma|    30.442 microns   | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|                                        |From new raw data
42|60 microns (IRAS)   | 5.111E-01 |+/-10  %|Jy                  |5.00E+12|  5.11E-01|+/-5.11E-02|Jy|1990IRASF.C...0000M|uncertainty| 60        microns   | Broad-band measurement|082757.9 +525527 (B1950)| Flux in fixed aperture|IRAS quality flag = 3                   |From new raw data
44|100 microns (IRAS)  | 9.511E-01 |+/-24  %|Jy                  |3.00E+12|  9.51E-01|+/-2.28E-01|Jy|1990IRASF.C...0000M|uncertainty| 100       microns   | Broad-band measurement|082757.9 +525527 (B1950)| Flux in fixed aperture|IRAS quality flag = 2                   |From new raw data
56|350 microns SHARC II| 386       |+/-32   |milliJy             |8.57E+11|  3.86E-01|+/-3.20E-02|Jy|2006ApJ...642..694B|1 sigma|     350   microns   | Broad-band measurement|08 31 41.70 +52 45 17.35 (J2000)| Flux integrated from map|                                        |From new raw data
58|450 microns SHARC II| 342       |+/-26   |milliJy             |6.66E+11|  3.42E-01|+/-2.60E-02|Jy|2006ApJ...642..694B|1 sigma|     450   microns   | Broad-band measurement|08 31 41.70 +52 45 17.35 (J2000)| Flux integrated from map|                                        |From new raw data
69|302 GHz (SMA)       | 60        |+/-12   | milliJy            |3.02E+11|  6.00E-02|+/-1.20E-02|Jy|2007ApJ...671L...5K|uncertainty|     302.4 GHz       | Broad-band measurement|| Flux integrated from map|                                        |From new raw data
70|250 GHz (PdBI)      | 34        |+/-0.55 |milliJy             |2.50E+11|  3.40E-02|+/-5.50E-04|Jy|2011ApJ...738L...6L|uncertainty|      250  GHz       | Broad-band measurement|| Flux integrated from map|                                        |From new raw data
71|245.905 GHz (IRAM)  | 31.4      |+/-2.0  |milliJy             |2.46E+11|  3.14E-02|+/-2.00E-03|Jy|2011ApJ...741L..38V|uncertainty|   245.905 GHz       | Broad-band measurement|| Flux integrated from map|                                        |From new raw data
72|236.797 GHz (PdBI)  | 26.6      |+/-1.3  |milliJy             |2.37E+11|  2.66E-02|+/-1.30E-03|Jy|2011ApJ...741L..38V|uncertainty|   236.797 GHz       | Broad-band measurement|| Flux integrated from map|                                        |From new raw data
74|201.166 GHz (IRAM)  | 16.5      |+/-0.8  |milliJy             |2.01E+11|  1.65E-02|+/-8.00E-04|Jy|2011ApJ...741L..38V|uncertainty|   201.166 GHz       | Broad-band measurement|| Flux integrated from map|                                        |From new raw data
75|153.132 GHz (PdBI)  | 5.4       |+/-0.3  |milliJy             |1.53E+11|  5.40E-03|+/-3.00E-04|Jy|2011ApJ...741L..38V|uncertainty|   153.132 GHz       | Broad-band measurement|| Flux integrated from map|                                        |From new raw data
78|110.7 GHz (CARMA)   | 2.17      |+/-0.19 |milliJy             |1.11E+11|  2.17E-03|+/-1.90E-04|Jy|2010ApJ...725.1032R|uncertainty|     110.7 GHz       | Broad-band measurement|| Flux integrated from map|                                        |From new raw data
79|108.6 GHz (CARMA)   | 2.08      |+/-0.22 |milliJy             |1.09E+11|  2.08E-03|+/-2.20E-04|Jy|2010ApJ...725.1032R|uncertainty|     108.6 GHz       | Broad-band measurement|| Flux integrated from map|                                        |From new raw data
80|105.4 GHz (CARMA)   | 2.04      |+/-0.08 |milliJy             |1.05E+11|  2.04E-03|+/-8.00E-05|Jy|2010ApJ...725.1032R|uncertainty|     105.4 GHz       | Broad-band measurement|| Flux integrated from map|                                        |From new raw data
82|90.8 GHz (PdBI)     | 1.2       |+/-0.13 |milliJy             |9.08E+10|  1.20E-03|+/-1.30E-04|Jy|2006ApJ...645L..17G|uncertainty| 90.797    GHz       | Broad-band measurement|08 31 41.73 +52 45 17.4 (J2000)| Flux integrated from map|Beam size = 1.46" x 1.20"               |From new raw data
83|87.0 GHz (GBT)      ||<0.1       | Jy                 |8.70E+10||1.00E-01|Jy|2004MNRAS.352..563C|1 sigma|      87.0 GHz       | Broad-band measurement|| Flux integrated from map|                                        |From new raw data
