
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-06-10T02:35:28PDT



Photometric Data for RGJ105209.31+572202.8 (z=2.112)

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|I (Cousins)             | 24.38     |+/-0.29 |mag                 |3.79E+14|  4.51E-07|+/-1.38E-07|Jy|2004ApJ...616...71S|1 sigma|    7900   A         | Broad-band measurement|| Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
2|K_s_ (2MASS)            | 20.24     |+/-0.30 |mag                 |1.38E+14|  5.35E-06|+/-1.70E-06|Jy|2004ApJ...616...71S|1 sigma|    2.17   microns   | Broad-band measurement|| Flux in fixed aperture|4" aperture                             |Averaged new and previously published data
3|24 microns (MIPS)       | 167.      |+/-47.0 |uJy             |1.27E+13|167.E-06|+/-47.E-06|Jy|2009ApJ...694.1517D|1rms uncertainty|     23.68 microns   | Broad-band measurement|12 37 11.89 +62 22 11.8 (J2000)| Flux integrated from map|                                        |From new raw data
4|70 microns (MIPS)       |           |<2.7    |mJy             |4.20E+12|        |2.7E-03|Jy|2009ApJ...699.1610H|3 sigma|     71.42 microns   | Broad-band measurement|221804.42 +002154.4 (J2000)| Flux in fixed aperture|                                        |From new raw data
5|350 microns (SHARC-II)  |           |<49.5   |mJy             |8.565E+11|      |49.5E-03|Jy|2005MNRAS.358..149P|3sigma uncertainty|     850   microns   | Broad-band measurement|12 37 11.7 +62 22 12 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
6|850 microns (SCUBA)     |           |<6.4    |milliJy            |3.53E+11|  |4.2E-03|Jy|2004ApJ...614..671C|3rms uncertainty|       850 microns   | Broad-band measurement|105209.31 +572202.8 (J2000)| Flux integrated from map|                                        |From new raw data
7|850 microns (SCUBA)     | 1.6       |+/-1.3  |milliJy            |3.53E+11|  1.60E-03|+/-1.30E-03|Jy|2004ApJ...614..671C|uncertainty|       850 microns   | Broad-band measurement|105209.31 +572202.8 (J2000)| Flux integrated from map|                                        |From new raw data
8|1200 microns (MAMBO)    |           |<2.7    |mJy             |2.50E+11|        |2.7E-03|Jy|2004MNRAS.354..779G|3 sigma uncertainty|      1200 microns   | Broad-band measurement|16 36 55.9 +40 59 12 (J2000)| Flux integrated from map|S/N = 3.66                              |From new raw data
9|1.4 GHz (VLA)           | 23        |+/-4    |microJy            |1.40E+09|  2.30E-05|+/-4.00E-06|Jy|2006MNRAS.371..963B|1 sigma|       1.4 GHz       | Broad-band measurement|10 52 09.450 +57 22 04.59 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
10|1.4 GHz (VLA)          | 34.5      |+/-5.5  |microJy            |1.40E+09|  34.5E-06|+/-5.5E-06|Jy|2006MNRAS.371..963B|1 sigma|       1.4 GHz       | Broad-band measurement|10 52 09.450 +57 22 04.59 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
