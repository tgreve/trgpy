

Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.


queryDateTime:2009-11-03T15:07:35PST






Photometric Data for MIPS16059 (z=2.326)

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|R (KPNO)            | 1.204     ||microJy             |4.66E+14|  1.20E-06||Jy|2007ApJ...658..778Y|no uncertainty reported|    6440   A         | Broad-band measurement|172428.44 +601533.2 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data
2|R (Cousins) m_aper  | 23.49     |+/-0.11 |mag                 |4.65E+14|  1.23E-06|+/-1.25E-07|Jy|2004AJ....128....1F|based on count statistics only|6440       A         | Broad-band measurement|172428.439 +601533.30 (J2000)| Flux in fixed aperture|3-arcsecond aperture                    |From new raw data
3|R (Cousins) m_aper  | 24.04     |+/-0.14 |mag                 |4.65E+14|  7.41E-07|+/-9.55E-08|Jy|2004AJ....128....1F|based on count statistics only|6440       A         | Broad-band measurement|172428.464 +601533.55 (J2000)| Flux in fixed aperture|3-arcsecond aperture                    |From new raw data
4|R (Cousins) m_tot   | 23.77     |+/-0.21 |mag                 |4.65E+14|  9.50E-07|+/-1.84E-07|Jy|2004AJ....128....1F|based on count statistics only|6440       A         | Broad-band measurement|172428.464 +601533.55 (J2000)| Total flux|                                        |From new raw data
5|R (Cousins) m_tot   | 23.47     |+/-0.12 |mag                 |4.65E+14|  1.25E-06|+/-1.38E-07|Jy|2004AJ....128....1F|based on count statistics only|6440       A         | Broad-band measurement|172428.439 +601533.30 (J2000)| Total flux|                                        |From new raw data
6|F160W (HST NICMOS)         | 20.29     ||mag                 |1.87E+14|  7.99E-06||Jy|2011ApJ...730..125Z|no uncertainty reported|      1.60 microns   | Broad-band measurement|| Flux integrated from map|                                        |From new raw data
7|F160W (HST NICMOS)         | 20.49     || mag                |1.86E+14|  6.65E-06||Jy|2008ApJ...680..232D|no uncertainty reported|      1.61 microns   | Broad-band measurement|17 24 28.34 +60 15 33.08 (J2000)| Flux integrated from map|                                        |From new raw data
8|3.6 microns (IRAC)  | 17        |+/-3    | microJy            |8.44E+13|  1.70E-05|+/-3.00E-06|Jy|2007ApJ...664..713S|uncertainty|   3.550   microns   | Broad-band measurement|| Flux in fixed aperture|7.3" diameter aperture                  |From reprocessed raw data
9|3.6 microns (IRAC)  ||<20.00     |microJy             |8.42E+13||2.00E-05|Jy|2005ApJS..161...41L|3sigma plate limit|3.56       microns   | Broad-band measurement|172428.34 +601533.1 (J2000)| Flux in fixed aperture|Aperture =       4.92 arcsec.           |From new raw data
10|4.5 microns (IRAC)  | 19        |+/-4    | microJy            |6.67E+13|  1.90E-05|+/-4.00E-06|Jy|2007ApJ...664..713S|uncertainty|   4.493   microns   | Broad-band measurement|| Flux in fixed aperture|7.3" diameter aperture                  |From reprocessed raw data
11|4.5 microns (IRAC)  ||<25.00     |microJy             |6.63E+13||2.50E-05|Jy|2005ApJS..161...41L|3sigma plate limit|4.52       microns   | Broad-band measurement|172428.34 +601533.1 (J2000)| Flux in fixed aperture|Aperture =       4.92 arcsec.           |From new raw data
12|5.8 microns (IRAC)  ||<100.00    |microJy             |5.23E+13||1.00E-04|Jy|2005ApJS..161...41L|3sigma plate limit|5.73       microns   | Broad-band measurement|172428.34 +601533.1 (J2000)| Flux in fixed aperture|Aperture =       4.92 arcsec.           |From new raw data
13|5.8 microns (IRAC)  | 33        |+/-14   | microJy            |5.23E+13|  3.30E-05|+/-1.40E-05|Jy|2007ApJ...664..713S|uncertainty|   5.731   microns   | Broad-band measurement|| Flux in fixed aperture|7.3" diameter aperture                  |From reprocessed raw data
16|8.0 microns (IRAC)  | 86.168    ||microJy             |3.81E+13|  8.62E-05||Jy|2007ApJ...658..778Y|no uncertainty reported|   7.872   microns   | Broad-band measurement|172428.44 +601533.2 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data
17|8.0 microns (IRAC)  | 66        |+/-15   | microJy            |3.81E+13|  6.60E-05|+/-1.50E-05|Jy|2007ApJ...664..713S|uncertainty|   7.872   microns   | Broad-band measurement|| Flux in fixed aperture|7.3" diameter aperture                  |From reprocessed raw data
18|8.0 microns (IRAC)  | 100.84    |+/-16.90|microJy             |3.79E+13|  1.01E-04|+/-1.69E-05|Jy|2005ApJS..161...41L|uncertainty|7.91       microns   | Broad-band measurement|172428.34 +601533.1 (J2000)| Flux in fixed aperture|Aperture =       4.92 arcsec.           |From new raw data
19|8 microns (IRAC) | 1.6       |+/-1   %|milliJy             |3.75E+13|  1.60E-03|+/-1.60E-05|Jy|2009ApJ...698.1682W|typical accuracy|         8 microns   | Broad-band measurement|17 24 28.44 +60 15 33.2 (J2000)| Peak flux|                                        |From reprocessed raw data
20|24 microns (MIPS)   | 1137.134  ||microJy             |1.27E+13|  1.14E-03||Jy|2007ApJ...658..778Y|no uncertainty reported|   23.68   microns   | Broad-band measurement|172428.44 +601533.2 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data; measurementmodified from published value
1|MIPS 24um           | 1.29     |+/-0.39 |milliJy             |1.27E+13|  1.29E-03|+/-0.39E-03 |Jy|1996AJ....111.1431B|uncertainty|1.49       GHz       | Broad-band measurement| | Peak flux|                                        |From new raw data
22|70 microns (MIPS)   | 6.2       |+/-2.4  | milliJy            |4.20E+12|  6.20E-03|+/-2.40E-03|Jy|2007ApJ...664..713S|estimated error|   71.42   microns   | Broad-band measurement|| Flux in fixed aperture|3 pixel radius aperture                 |From reprocessed raw data
2|MIPS 70um           |          |<7.2    |milliJy             |4.20E+12|          |7.2E-03|Jy|2010Natur.464..733S|3sigma uncertainty|     71.42 microns   | Broad-band measurement|21 35 11.6 -01 02 52.0 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
3|MIPS 160um          |          |<30     |milliJy             |1.92E+12|          |30.0E-03|Jy|2009A&A...502..541E|3 sigma|     155.9 microns   | Broad-band measurement| | Flux in fixed aperture|                                        |From reprocessed raw data
4|MAMBO 1200um        | 1.20     |+/-0.66 |milliJy             |2.50E+11|  1.20E-03|+/-0.66E-03|Jy|2004MNRAS.354..779G|uncertainty|      1200 microns   | Broad-band measurement|16 37 06.7 +40 53 15 (J2000)| Flux integrated from map|S/N = 3.81                              |From new raw data
5|VLA 1.4GHz          | 0.57     |+/-0.03 |milliJy             |1.4E9   |  0.57E-3 |+/-0.03E-3|Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
