
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-02-19T12:35:26PST



Photometric Data for ERO J164502+4626.4

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|4400 Angstroms      | 0.16      |+/-0.07 |microJy             |6.81E+14|  1.60E-07|+/-7.00E-08|Jy|1999ApJ...519..610D|uncertainty| 4400      Angstroms | Broad-band measurement|164502.36 +462625.5 (J2000)| Flux in fixed aperture|3" aperture                             |From reprocessed raw data
2|R_aper (WHT) AB     | 25.189    | |mag                 |4.70E+14|  3.05E-07| |Jy|2005MNRAS.360..685C|no uncertainty reported|    6380   A         | Broad-band measurement|16 45 02.30 +46 26 26.23 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data; derived from a fluxin a different band and a color
3|7930 Angstroms      | 0.52      |+/-0.06 |microJy             |3.78E+14|  5.20E-07|+/-6.00E-08|Jy|1999ApJ...519..610D|uncertainty| 7924      Angstroms | Broad-band measurement|164502.36 +462625.5 (J2000)| Flux in fixed aperture|3" aperture                             |From new raw data
4|1.2 microns         | 6.4       |+/-2.1  |microJy             |2.40E+14|  6.40E-06|+/-2.10E-06|Jy|1999ApJ...519..610D|uncertainty| 1.2       microns   | Broad-band measurement|164502.36 +462625.5 (J2000)| Flux in fixed aperture|3" aperture                             |From reprocessed raw data; Standard Caltech JHKL filtersassumed
5|1.6 microns         | 14.8      |+/-3.6  |microJy             |1.82E+14|  1.48E-05|+/-3.60E-06|Jy|1999ApJ...519..610D|uncertainty| 1.6       microns   | Broad-band measurement|164502.36 +462625.5 (J2000)| Flux in fixed aperture|3" aperture                             |Averaged from previously published data; Standard CaltechJHKL filters assumed
6|K_aper (UKIRT) AB   | 20.44     | |mag                 |1.37E+14|  2.42E-05| |Jy|2005MNRAS.360..685C|no uncertainty reported|   2.195   microns   | Broad-band measurement|16 45 02.30 +46 26 26.23 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
7|2.2 microns         | 27.7      |+/-0.6  |microJy             |1.36E+14|  2.77E-05|+/-6.00E-07|Jy|1999ApJ...519..610D|uncertainty| 2.2       microns   | Broad-band measurement|164502.36 +462625.5 (J2000)| Flux in fixed aperture|3" aperture                             |Averaged from previously published data; Standard CaltechJHKL filters assumed
8|IRAS 12 microns     | |<75        |milliJy             |2.50E+13| |7.50E-02|Jy|1999ApJ...519..610D|3sisgma uncertainty reported| 12        microns   | Broad-band measurement|164502.36 +462625.5 (J2000)| Integrated from scans|                                        |Averaged from previously published data
9|IRAS 25 microns     | |<60        |milliJy             |1.20E+13| |6.00E-02|Jy|1999ApJ...519..610D|3sisgma uncertainty reported| 25        microns   | Broad-band measurement|164502.36 +462625.5 (J2000)| Integrated from scans|                                        |Averaged from previously published data
10|IRAS 60 microns     | |<84        |milliJy             |5.00E+12| |8.40E-02|Jy|1999ApJ...519..610D|3sisgma uncertainty reported| 60        microns   | Broad-band measurement|164502.36 +462625.5 (J2000)| Integrated from scans|                                        |Averaged from previously published data
11|IRAS 100 microns    | |<270       |milliJy             |3.00E+12| |2.70E-01|Jy|1999ApJ...519..610D|3sisgma uncertainty reported| 100       microns   | Broad-band measurement|164502.36 +462625.5 (J2000)| Integrated from scans|                                        |Averaged from previously published data
12|SCUBA 450 microns   | 32.3      |+/-8.5  |milliJy             |6.66E+11|  3.23E-02|+/-8.50E-03|Jy|1999ApJ...519..610D|uncertainty| 450       microns   | Broad-band measurement|164502.36 +462625.5 (J2000)| Flux integrated from map|                                        |From new raw data
13|SCUBA 850 microns   | 4.89      |+/-0.74 |milliJy             |3.53E+11|  4.89E-03|+/-7.40E-04|Jy|1999ApJ...519..610D|uncertainty| 850       microns   | Broad-band measurement|164502.36 +462625.5 (J2000)| Flux integrated from map|                                        |From new raw data
14|SCUBA 1350 microns  | 2.13      |+/-0.63 |milliJy             |2.22E+11|  2.13E-03|+/-6.30E-04|Jy|1999ApJ...519..610D|uncertainty| 1350      microns   | Broad-band measurement|164502.36 +462625.5 (J2000)| Flux integrated from map|                                        |From new raw data
15|VLA 3.6 cm          | 35        |+/-11   |microJy             |8.33E+09|  3.50E-05|+/-1.10E-05|Jy|1999ApJ...519..610D|uncertainty| 3.6       cm        | Broad-band measurement|164502.36 +462625.5 (J2000)| Flux integrated from map|                                        |From new raw data
16|VLA 20 cm           | |<300       |microJy             |1.50E+09| |3.00E-04|Jy|1999ApJ...519..610D|3sigma uncertainty reported| 20        cm        | Broad-band measurement|164502.36 +462625.5 (J2000)| Not reported in paper|                                        |Averaged from previously published data
