
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-07-10T12:59:00PDT



Photometric Data for LEDA 2830749

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|J_s (VLT)           | 4.1       |+/-1.5  |microJy             |2.50E+14|  4.10E-06|+/-1.50E-06|Jy|2006MNRAS.366L...1V|uncertainty|     1.2   microns   | Broad-band measurement|| Corrected to total flux from single aperture measurement|Flux corrected for line emission        |From new raw data
2|F160W (HST/NIC)     | 1.7       |+/-1.2  |microJy             |1.87E+14|  1.70E-06|+/-1.20E-06|Jy|2006MNRAS.366L...1V|uncertainty|     1.6   microns   | Broad-band measurement|| Corrected to total flux from single aperture measurement|Flux corrected for line emission        |From new raw data
3|K_s (VLT)           | 4.8       |+/-1.8  |microJy             |1.36E+14|  4.80E-06|+/-1.80E-06|Jy|2006MNRAS.366L...1V|uncertainty|     2.2   microns   | Broad-band measurement|| Corrected to total flux from single aperture measurement|Flux corrected for line emission        |From new raw data
4|3.6 microns (IRAC)  | 28.1      |+/-3.3  | microJy            |8.44E+13|  2.81E-05|+/-3.30E-06|Jy|2007ApJS..171..353S|uncertainty|   3.550   microns   | Broad-band measurement|21 06 58.1 -24 05 11.00 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
5|3.6 microns (IRAC)  | 27        |+/-3    |microJy             |8.33E+13|  2.70E-05|+/-3.00E-06|Jy|2006MNRAS.366L...1V|uncertainty|     3.6   microns   | Broad-band measurement|| Corrected to total flux from single aperture measurement|                                        |From new raw data
6|4.5 microns (IRAC)  | 29.7      |+/-3.5  | microJy            |6.67E+13|  2.97E-05|+/-3.50E-06|Jy|2007ApJS..171..353S|uncertainty|   4.493   microns   | Broad-band measurement|21 06 58.1 -24 05 11.00 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
7|4.5 microns (IRAC)  | 29        |+/-3    |microJy             |6.66E+13|  2.90E-05|+/-3.00E-06|Jy|2006MNRAS.366L...1V|uncertainty|     4.5   microns   | Broad-band measurement|| Corrected to total flux from single aperture measurement|                                        |From new raw data
8|5.8 microns (IRAC)  | 32        |+/-7    |microJy             |5.26E+13|  3.20E-05|+/-7.00E-06|Jy|2006MNRAS.366L...1V|uncertainty|     5.7   microns   | Broad-band measurement|| Corrected to total flux from single aperture measurement|                                        |From new raw data
9|5.8 microns (IRAC)  | 32.8      |+/-10.0 | microJy            |5.23E+13|  3.28E-05|+/-1.00E-05|Jy|2007ApJS..171..353S|uncertainty|   5.731   microns   | Broad-band measurement|21 06 58.1 -24 05 11.00 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
10|8.0 microns (IRAC)  ||<36.3      | microJy            |3.81E+13||3.63E-05|Jy|2007ApJS..171..353S|3 sigma|   7.872   microns   | Broad-band measurement|21 06 58.1 -24 05 11.00 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data
11|8.0 microns (IRAC)  ||<35        |microJy             |3.75E+13||3.50E-05|Jy|2006MNRAS.366L...1V|no uncertainty reported|     8.0   microns   | Broad-band measurement|| Corrected to total flux from single aperture measurement|                                        |From new raw data
12|16.0 microns (IRS)  | 72        |+/-18   |microJy             |1.87E+13|  7.20E-05|+/-1.80E-05|Jy|2006MNRAS.366L...1V|uncertainty|    16.0   microns   | Broad-band measurement|| Corrected to total flux from single aperture measurement|                                        |From new raw data
13|16 microns (IRS)    | 121.0     |+/-47.0 | microJy            |1.87E+13|  1.21E-04|+/-4.70E-05|Jy|2007ApJS..171..353S|uncertainty|      16   microns   | Broad-band measurement|21 06 58.1 -24 05 11.00 (J2000)| Flux in fixed aperture|6" diameter aperture                    |From reprocessed raw data
14|4.85 GHz            | 107       |+/-12   |milliJy             |4.85E+09|  1.07E-01|+/-1.20E-02|Jy|1994ApJS...90..179G|rms noise|4.85       GHz       | Broad-band measurement|210658.3 -240444 (J2000)| Modelled datum|                                        |From new raw data; Corrected for contaminating sources
15|408 MHz             | 1.80      |+/-0.09 |Jy                  |4.08E+08|  1.80E+00|+/-9.00E-02|Jy|1981MNRAS.194..693L|rms noise|408        MHz       | Broad-band measurement|210404.6 -241723 (B1950)| Modelled datum|                                        |From new raw data; Corrected for contaminating sources
16|365 MHz (Texas)     | 2.232     |+/-0.120|Jy                  |3.65E+08|  2.23E+00|+/-1.20E-01|Jy|1996AJ....111.1945D|internal error|365        MHz       | Broad-band measurement; obtained by interpolation over frequency|210403.980 -241711.79 (B1950)| Integrated from scans|Model:D;MFlag:+;EFlag:+;LFlag:+.        |From new raw data
17|74 MHz (VLA)        | 10.51     |+/-1.15 | Jy                 |7.38E+07|  1.05E+01|+/-1.15E+00|Jy|2007AJ....134.1245C|rms uncertainty|      73.8 MHz       | Broad-band measurement|21 06 58.10 -24 05 08.7 (J2000)| Flux integrated from map|Corrected for clean bias                |From new raw data
