


Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.





Photometric Data GN20.2a, z=4.05

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|R (Keck II) AB       | 25.44    | | mag       |4.62E+14|  2.42E-07| |Jy|2004AJ....127.3121W|no uncertainty reported|   648.7   A         | Broad-band measurement|12 37 11.815 +62 22 11.84 (J2000)| Total flux|           
2|i (775HST) AB        | 24.7     | | mag       |3.897E+14|  4.78E-07| |Jy|2004AJ....127.3121W|no uncertainty reported|   648.7   A         | Broad-band measurement|12 37 11.815 +62 22 11.84 (J2000)| Total flux|           
3|3.6 microns IRAC     | 3.87     |+/-0.55|uJy  |8.44E+13|  3.87E-06|+/-0.55E-06|Jy|2005ApJ...635..853B|uncertainty|   3.550   microns   | Broad-band measurement|123707.21 +621408.1 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged new and previously published data
4|4.5um (Spitzer)      | 4.1      |+/-0.4 |uJy  | 6.67E13 | 4.1E-6  |+/-0.4E-6 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
5|4.5um (Spitzer)      | 3.89     |+/-0.51|uJy  | 6.67E13 | 3.89E-6  |+/-0.51E-6 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
6|5.7 microns (IRAC)   | 6.06     |+/-0.98|uJy  |5.23E+13|  6.06E-06|+/-0.98E-06|Jy|2008ApJ...675..262R|uncertainty|     5.731 microns   | Broad-band measurement|14 01 04.96 +02 52 24.8 (J2000)| Flux in fixed aperture|                                        |From new raw data
7|8.0um (Spitzer)      | 9.8      |+/-1.0 |uJy  | 3.75E13 | 9.8E-6  |+/-1.0E-6 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
9|8.0um (Spitzer)      | 9.36     |+/-1.14|uJy  | 3.75E13 | 9.36E-6  |+/-1.14E-6 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
10|24um (Spitzer)      | 30.2     |+/-5.6 |uJy  | 1.25E13 | 30.2E-6 |+/-5.6E-6 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
11|850um (SCUBA)       | 9.9      |+/-2.3 |mJy  | 3.529E11| 9.9E-3  |+/-2.3E-3 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
12|2mm (PdBI)          | 0.7      |+/-0.2 |mJy  | 136.96E9| 0.7E-03|+/-0.2E-03 |Jy |2003MNRAS.343..293M|rms uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
13|3.3mm (IRAM)        |          |<0.20  |mJy  | 9.09E10 | |0.20E-03     |Jy |2003MNRAS.343..293M|3rms uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
14|1.4GHz (VLA)        | 180.7    |+/-8.4 |uJy  | 1.4E9   | 180.7E-6|+/-8.4E-6 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
