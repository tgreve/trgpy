
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-06-11T21:22:18PDT



Photometric Data for GOODS J123707.21+621408.1

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|1.4 GHz (VLA)       | 30.      |+/-8.  | microJy            |1.40E+09|  39.E-06|+/-8.E-06|Jy|2007MNRAS.380..199I|rms uncertainty|       1.4 GHz       | Broad-band measurement|10 52 28.995 +57 22 22.42 (J2000)| Flux integrated from map|                                        |From reprocessed raw data
