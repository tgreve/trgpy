
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-06-16T05:44:23PDT



Photometric Data for SDSS J141859.16+524716.5

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|FUV (GALEX) AB      ||>24.0262   |mag                 |1.95E+15||8.90E-07|Jy|2012GMSC..C...0000S|3 sigma|1538.6     A         | Broad-band measurement|214.74631440188 52.787906788771 (J2000)| Flux integrated from map|upper limit inside NUV Kron aperture    |From new raw data
2|FUV (GALEX) AB      | 25.3997   |+/-0.586945|mag                 |1.95E+15|  2.51E-07|+/-1.36E-07|Jy|2012GMSC..C...0000S|uncertainty|1538.6     A         | Broad-band measurement|214.74631440188 52.787906788771 (J2000)| Flux in fixed aperture|Flux in 7.5 arcsec diameter aperture    |From new raw data
3|NUV (GALEX) AB      | 23.7387   |+/-0.212787|mag                 |1.29E+15|  1.16E-06|+/-2.27E-07|Jy|2012GMSC..C...0000S|uncertainty|2315.7     A         | Broad-band measurement|214.74631440188 52.787906788771 (J2000)| Flux integrated from map|Kron flux in elliptical aperture        |From new raw data
4|NUV (GALEX) AB      | 23.9732   |+/-0.132455|mag                 |1.29E+15|  9.35E-07|+/-1.14E-07|Jy|2012GMSC..C...0000S|uncertainty|2315.7     A         | Broad-band measurement|214.74631440188 52.787906788771 (J2000)| Flux in fixed aperture|Flux in 7.5 arcsec diameter aperture    |From new raw data
5|u (SDSS CModel) AB  | 22.095    ||asinh mag           |8.36E+14|  5.42E-06||Jy|2007SDSS6.C...0000:|no uncertainty reported|3585       A         | Broad-band measurement|214.7465123314 52.7879206934 (J2000)| Modelled datum|SDSS flags: CANONICAL_CENTER - used canonical, not local, center; NOPETRO - no Petrosian radius could be determined; BAD_RADIAL - some low S/N radial points; PETROFAINT - Petrosian radius measured at very low surface brightness; ELLIPFAINT - no isophotal fits performed; AMOMENT_FAINT - too faint for adaptive moments;|From new raw data
6|u (SDSS Model) AB   | 23.039    |+/-0.603|asinh mag           |8.36E+14|  2.17E-06|+/-1.34E-06|Jy|2007SDSS6.C...0000:|based on count statistics only|3585       A         | Broad-band measurement|214.7465123314 52.7879206934 (J2000)| Modelled datum|SDSS flags: CANONICAL_CENTER - used canonical, not local, center; NOPETRO - no Petrosian radius could be determined; BAD_RADIAL - some low S/N radial points; PETROFAINT - Petrosian radius measured at very low surface brightness; ELLIPFAINT - no isophotal fits performed; AMOMENT_FAINT - too faint for adaptive moments;|From new raw data
7|u (SDSS PSF) AB     | 23.276    |+/-0.475|asinh mag           |8.36E+14|  1.69E-06|+/-8.72E-07|Jy|2007SDSS6.C...0000:|based on count statistics only|3585       A         | Broad-band measurement|214.7465123314 52.7879206934 (J2000)| Modelled datum|SDSS flags: CANONICAL_CENTER - used canonical, not local, center; NOPETRO - no Petrosian radius could be determined; BAD_RADIAL - some low S/N radial points; PETROFAINT - Petrosian radius measured at very low surface brightness; ELLIPFAINT - no isophotal fits performed; AMOMENT_FAINT - too faint for adaptive moments;|From new raw data
8|g (SDSS Model) AB   | 22.136    |+/-0.148|asinh mag           |6.17E+14|  5.06E-06|+/-6.95E-07|Jy|2007SDSS6.C...0000:|based on count statistics only|4858       A         | Broad-band measurement|214.7465123314 52.7879206934 (J2000)| Modelled datum|SDSS flags: NOPETRO - no Petrosian radius could be determined; BAD_RADIAL - some low S/N radial points; PETROFAINT - Petrosian radius measured at very low surface brightness; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
9|g (SDSS CModel) AB  | 22.181    ||asinh mag           |6.17E+14|  4.85E-06||Jy|2007SDSS6.C...0000:|no uncertainty reported|4858       A         | Broad-band measurement|214.7465123314 52.7879206934 (J2000)| Modelled datum|SDSS flags: NOPETRO - no Petrosian radius could be determined; BAD_RADIAL - some low S/N radial points; PETROFAINT - Petrosian radius measured at very low surface brightness; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
10|g (SDSS PSF) AB     | 22.739    |+/-0.158|asinh mag           |6.17E+14|  2.88E-06|+/-4.29E-07|Jy|2007SDSS6.C...0000:|based on count statistics only|4858       A         | Broad-band measurement|214.7465123314 52.7879206934 (J2000)| Modelled datum|SDSS flags: NOPETRO - no Petrosian radius could be determined; BAD_RADIAL - some low S/N radial points; PETROFAINT - Petrosian radius measured at very low surface brightness; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
11|r (SDSS CModel) AB  | 21.648    ||asinh mag           |4.77E+14|  7.93E-06||Jy|2007SDSS6.C...0000:|no uncertainty reported|6290       A         | Broad-band measurement|214.7465123314 52.7879206934 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding; CANONICAL_BAND - this band was primary (usually r);|From new raw data
12|r (SDSS Model) AB   | 21.647    |+/-0.112|asinh mag           |4.77E+14|  7.94E-06|+/-8.24E-07|Jy|2007SDSS6.C...0000:|based on count statistics only|6290       A         | Broad-band measurement|214.7465123314 52.7879206934 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding; CANONICAL_BAND - this band was primary (usually r);|From new raw data
13|r (SDSS PSF) AB     | 22.218    |+/-0.116|asinh mag           |4.77E+14|  4.67E-06|+/-5.07E-07|Jy|2007SDSS6.C...0000:|based on count statistics only|6290       A         | Broad-band measurement|214.7465123314 52.7879206934 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding; CANONICAL_BAND - this band was primary (usually r);|From new raw data
14|i (SDSS Model) AB   | 21.581    |+/-0.160|asinh mag           |3.89E+14|  8.41E-06|+/-1.25E-06|Jy|2007SDSS6.C...0000:|based on count statistics only|7706       A         | Broad-band measurement|214.7465123314 52.7879206934 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
15|i (SDSS CModel) AB  | 21.662    ||asinh mag           |3.89E+14|  7.80E-06||Jy|2007SDSS6.C...0000:|no uncertainty reported|7706       A         | Broad-band measurement|214.7465123314 52.7879206934 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
16|i (SDSS PSF) AB     | 22.017    |+/-0.144|asinh mag           |3.89E+14|  5.59E-06|+/-7.61E-07|Jy|2007SDSS6.C...0000:|based on count statistics only|7706       A         | Broad-band measurement|214.7465123314 52.7879206934 (J2000)| Modelled datum|SDSS flags: BAD_RADIAL - some low S/N radial points; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
17|z (SDSS Model) AB   | 20.472    |+/-0.206|asinh mag           |3.25E+14|  2.28E-05|+/-4.44E-06|Jy|2007SDSS6.C...0000:|based on count statistics only|9222       A         | Broad-band measurement|214.7465123314 52.7879206934 (J2000)| Modelled datum|SDSS flags: MANYPETRO - more than one Petrosian radius; BAD_RADIAL - some low S/N radial points; ELLIPFAINT - no isophotal fits performed; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
18|z (SDSS PSF) AB     | 20.873    |+/-0.184|asinh mag           |3.25E+14|  1.55E-05|+/-2.78E-06|Jy|2007SDSS6.C...0000:|based on count statistics only|9222       A         | Broad-band measurement|214.7465123314 52.7879206934 (J2000)| Modelled datum|SDSS flags: MANYPETRO - more than one Petrosian radius; BAD_RADIAL - some low S/N radial points; ELLIPFAINT - no isophotal fits performed; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
19|z (SDSS CModel) AB  | 19.884    ||asinh mag           |3.25E+14|  3.95E-05||Jy|2007SDSS6.C...0000:|no uncertainty reported|9222       A         | Broad-band measurement|214.7465123314 52.7879206934 (J2000)| Modelled datum|SDSS flags: MANYPETRO - more than one Petrosian radius; BAD_RADIAL - some low S/N radial points; ELLIPFAINT - no isophotal fits performed; BINNED1 - detected at >=5 sigma in original imaging frame; BINNED_CENTER - image was binned while centroiding;|From new raw data
