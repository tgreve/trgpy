
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-07-08T05:13:01PDT



Photometric Data for GOODS J123712.15+621754.3

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|4.0-8 keV (Chandra) | 0.70E-15  ||ergs cm^-2^ s^-1^   |1.45E+18|  4.82E-11||Jy|2003AJ....126..539A|no uncertainty reported|       6   keV       | Broad-band measurement|12 37 12.12 +62 17 53.9 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
2|4-8 keV (Chandra)   ||<0.61E-15  |erg cm^-2^ s^-1^    |1.45E+18||4.21E-11|Jy|2001AJ....122.2810B|no uncertainty reported|       6   keV       | Broad-band measurement|12 37 12.12 +62 17 53.9 (J2000)| Flux in fixed aperture|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
3|2-8 keV (Chandra)   | 1.12E-15  |+/-4   %|erg cm^-2^ s^-1^    |1.21E+18|  9.26E-11|+/-3.70E-12|Jy|2001AJ....122.2810B|estimated error|       5   keV       | Broad-band measurement|12 37 12.12 +62 17 53.9 (J2000)| Flux in fixed aperture|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
4|2.0-8 keV (Chandra) | 1.14E-15  ||ergs cm^-2^ s^-1^   |1.21E+18|  9.43E-11||Jy|2003AJ....126..539A|no uncertainty reported|       5   keV       | Broad-band measurement|12 37 12.12 +62 17 53.9 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
5|0.5-8 keV (Chandra) | 1.93E-15  |+/-4   %|erg cm^-2^ s^-1^    |1.03E+18|  1.87E-10|+/-7.50E-12|Jy|2001AJ....122.2810B|estimated error|    4.25   keV       | Broad-band measurement|12 37 12.12 +62 17 53.9 (J2000)| Flux in fixed aperture|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
6|0.5-8 keV (Chandra) | 1.95E-15  ||ergs cm^-2^ s^-1^   |1.03E+18|  1.90E-10||Jy|2003AJ....126..539A|no uncertainty reported|    4.25   keV       | Broad-band measurement|12 37 12.12 +62 17 53.9 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
7|2.0-4 keV (Chandra) | 0.51E-15  ||ergs cm^-2^ s^-1^   |7.25E+17|  7.03E-11||Jy|2003AJ....126..539A|no uncertainty reported|       3   keV       | Broad-band measurement|12 37 12.12 +62 17 53.9 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
8|1.0-2 keV (Chandra) | 0.47E-15  ||ergs cm^-2^ s^-1^   |3.63E+17|  1.30E-10||Jy|2003AJ....126..539A|no uncertainty reported|     1.5   keV       | Broad-band measurement|12 37 12.12 +62 17 53.9 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
9|0.5-2 keV (Chandra) | 0.78E-15  ||ergs cm^-2^ s^-1^   |3.02E+17|  2.58E-10||Jy|2003AJ....126..539A|no uncertainty reported|    1.25   keV       | Broad-band measurement|12 37 12.12 +62 17 53.9 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
10|0.5-2 keV (Chandra) | 0.84E-15  |+/-4   %|erg cm^-2^ s^-1^    |3.02E+17|  2.78E-10|+/-1.11E-11|Jy|2001AJ....122.2810B|estimated error|    1.25   keV       | Broad-band measurement|12 37 12.12 +62 17 53.9 (J2000)| Flux in fixed aperture|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
11|0.5-1 keV (Chandra) | 0.36E-15  ||ergs cm^-2^ s^-1^   |1.81E+17|  1.98E-10||Jy|2003AJ....126..539A|no uncertainty reported|    0.75   keV       | Broad-band measurement|12 37 12.12 +62 17 53.9 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
12|U (KPNO) AB         | 25.3      || mag                |8.22E+14|  2.75E-07||Jy|2004AJ....127.3137C|no uncertainty reported| 3647.65   A         | Broad-band measurement|189.300629 +62.29843 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
13|F435W (HST/ACS) AB      | 22.683    |+/-0.014|mag                 |6.92E+14|  3.07E-06|+/-3.96E-08|Jy|2011ApJ...734..121S|uncertainty|      4333 A         | Broad-band measurement|189.300629 62.298428 (J2000)| Total flux|                                        |From reprocessed raw data
14|F435W (HST/ACS) AB      | 22.84     |+/-0.18 |mag                 |6.92E+14|  2.65E-06|+/-4.40E-07|Jy|2011ApJ...734..121S|uncertainty|      4333 A         | Broad-band measurement|189.300629 62.298428 (J2000)| Modelled datum|Host galaxy mag                         |From reprocessed raw data
15|F435W (HST/ACS) AB      | 24.89     |+/-0.14 |mag                 |6.92E+14|  4.02E-07|+/-5.18E-08|Jy|2011ApJ...734..121S|uncertainty|      4333 A         | Broad-band measurement|189.300629 62.298428 (J2000)| Modelled datum|Central point source mag                |From reprocessed raw data
16|B (Subaru) AB       | 25.3      || mag                |6.77E+14|  2.75E-07||Jy|2004AJ....127.3137C|no uncertainty reported| 4427.60   A         | Broad-band measurement|189.300629 +62.29843 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
17|V (Subaru) AB       | 24.7      || mag                |5.48E+14|  4.79E-07||Jy|2004AJ....127.3137C|no uncertainty reported| 5471.22   A         | Broad-band measurement|189.300629 +62.29843 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
18|R (Keck II) AB      | 24.39     || mag                |4.62E+14|  6.37E-07||Jy|2004AJ....127.3121W|no uncertainty reported|   648.7   A         | Broad-band measurement|12 37 12.130 +62 17 54.16 (J2000)| Total flux|                                        |From new raw data
19|R (Subaru) AB       | 24.0      || mag                |4.59E+14|  9.12E-07||Jy|2004AJ....127.3137C|no uncertainty reported| 6534.16   A         | Broad-band measurement|189.300629 +62.29843 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
20|R (Subaru) AB       | 24.02     ||mag                 |4.58E+14|  8.95E-07||Jy|2007MNRAS.377..203G|no uncertainty reported|    6550   A         | Broad-band measurement|12 37 12.12 +62 17 53.9 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
21|I (Subaru) AB       | 23.4      || mag                |3.76E+14|  1.59E-06||Jy|2004AJ....127.3137C|no uncertainty reported| 7975.89   A         | Broad-band measurement|189.300629 +62.29843 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
22|z' (Subaru) AB      | 22.8      || mag                |3.31E+14|  2.75E-06||Jy|2004AJ....127.3137C|no uncertainty reported| 9069.21   A         | Broad-band measurement|189.300629 +62.29843 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
23|HK' (UH) AB         | 21.0      || mag                |1.58E+14|  1.45E-05||Jy|2004AJ....127.3137C|no uncertainty reported|18947.38   A         | Broad-band measurement|189.300629 +62.29843 (J2000)| Corrected to total flux from single aperture measurement|                                        |Averaged from previously published data
24|3.6 microns (IRAC)  | 34.40     |+/-1.72 |microJy             |8.44E+13|  3.44E-05|+/-1.72E-06|Jy|2011AJ....141....1T|rms uncertainty|     3.550 microns   | Broad-band measurement|189.300690 62.298355 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
25|3.6 microns (IRAC)  | 34.40     |+/-0.05 |microJy             |8.44E+13|  3.44E-05|+/-5.00E-08|Jy|2007MNRAS.377..203G|uncertainty|   3.550   microns   | Broad-band measurement|12 37 12.12 +62 17 53.9 (J2000)| Corrected to total flux from single aperture measurement|                                        |From reprocessed raw data
26|4.5 microns (IRAC)  | 33.30     |+/-1.67 |microJy             |6.67E+13|  3.33E-05|+/-1.67E-06|Jy|2011AJ....141....1T|rms uncertainty|     4.493 microns   | Broad-band measurement|189.300690 62.298355 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
27|4.5 microns (IRAC)  | 34.15     |+/-0.09 |microJy             |6.67E+13|  3.42E-05|+/-9.00E-08|Jy|2007MNRAS.377..203G|uncertainty|   4.493   microns   | Broad-band measurement|12 37 12.12 +62 17 53.9 (J2000)| Corrected to total flux from single aperture measurement|                                        |From reprocessed raw data
28|5.8 microns (IRAC)  | 25.50     |+/-1.34 |microJy             |5.23E+13|  2.55E-05|+/-1.34E-06|Jy|2011AJ....141....1T|rms uncertainty|     5.731 microns   | Broad-band measurement|189.300690 62.298355 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
29|5.8 microns (IRAC)  | 25.79     |+/-0.44 |microJy             |5.23E+13|  2.58E-05|+/-4.40E-07|Jy|2007MNRAS.377..203G|uncertainty|   5.731   microns   | Broad-band measurement|12 37 12.12 +62 17 53.9 (J2000)| Corrected to total flux from single aperture measurement|                                        |From reprocessed raw data
30|8.0 microns (IRAC)  | 29.68     |+/-0.46 |microJy             |3.81E+13|  2.97E-05|+/-4.60E-07|Jy|2007MNRAS.377..203G|uncertainty|   7.872   microns   | Broad-band measurement|12 37 12.12 +62 17 53.9 (J2000)| Corrected to total flux from single aperture measurement|                                        |From reprocessed raw data
31|8.0 microns (IRAC)  | 29.50     |+/-1.55 |microJy             |3.81E+13|  2.95E-05|+/-1.55E-06|Jy|2011AJ....141....1T|rms uncertainty|     7.872 microns   | Broad-band measurement|189.300690 62.298355 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
32|16 microns (IRS)    | 183.8     |+/-10.5 |microJy             |1.90E+13|  1.84E-04|+/-1.05E-05|Jy|2011AJ....141....1T|rms uncertainty|      15.8 microns   | Broad-band measurement|189.300690 62.298355 (J2000)| From fitting to map|                                        |From new raw data
33|24 microns (MIPS)   | 139.56    |+/-5.01 |microJy             |1.27E+13|  1.40E-04|+/-5.01E-06|Jy|2007MNRAS.377..203G|uncertainty|   23.68   microns   | Broad-band measurement|12 37 12.12 +62 17 53.9 (J2000)| Corrected to total flux from single aperture measurement|                                        |From reprocessed raw data
34|24 microns (MIPS)   | 144.0     |+/-3.8  |microJy             |1.27E+13|  1.44E-04|+/-3.80E-06|Jy|2011AJ....141....1T|rms uncertainty|     23.68 microns   | Broad-band measurement|189.300690 62.298355 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
35|24 microns (MIPS)   | 154.6     |+/-2.6  |microJy             |1.27E+13|  1.55E-04|+/-2.60E-06|Jy|2011A&A...528A..35M|uncertainty|     23.68 microns   | Broad-band measurement|12 37 12.17 +62 17 54.01 (J2000)| Flux integrated from map|                                        |From new raw data
1|MIPS 24 microns      | 153.    |+/-5.0 |microJy         |1.25E+13 |  153.E-06|+/-5.0E-06  |Jy |1990IRASF.C...0000M|3sigma uncertainty| 25        microns   | Broad-band measurement|115813.1 +302058 (B1950)| Flux in fixed aperture|                                        |From new raw data
36|70 microns (MIPS)   ||<2.1       |milliJy             |4.20E+12||2.10E-03|Jy|2011A&A...528A..35M|no uncertainty reported|     71.42 microns   | Broad-band measurement|12 37 12.17 +62 17 54.01 (J2000)| Flux integrated from map|                                        |From new raw data
2|70 microns (PACS)    |         |<2.0   |mJy             |4.283e+12|          |2.0E-03     |Jy |2.40e+01           |3sigma   |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
3|100 microns (PACS)   | 2.6     |+/-0.3 |mJy             |2.998e+12|  2.6E-03 |+/-0.3E-03  |Jy |2.40e+01           |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
4|160 microns (PACS)   | 3.5     |+/-0.7 |mJy             |1.874e+12|  3.5E-03 |+/-0.7E-03  |Jy |2.40e+01           |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
5|250 microns (SPIRE)  | 6.2     |+/-2.5 |mJy             |1.199e+12|  6.2E-03 |+/-2.5e-03  |Jy |2.40e+01           |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
6|350 microns (SPIRE)  |         |<9.0   |mJy             |8.565e+11|          |9.0e-03     |Jy |2.40e+01           |3sigma   |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
7|500 microns (SPIRE)  |         |<12.0  |mJy             |5.996e+11|          |12.0e-03    |Jy |2.40e+01           |3sigma   |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
8|1160 microns (Penner)|         |<1.7   |mJy             |2.58442E+11|        |1.7E-03     |Jy |2004MNRAS.354..779G|3sigma uncertainty|      1200 microns   | Broad-band measurement|16 36 55.9 +40 59 12 (J2000)| Flux integrated from map|S/N = 3.66                              |From new raw data
