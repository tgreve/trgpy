
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-05-28T01:42:09PDT



Photometric Data for PEPJ123615+621008 (z=1.027)

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|2-8 keV (Chandra)   ||<-15.53    |log(erg/cm^2^/s)    |1.21E+18||2.44E-11|Jy|2008ApJ...681.1163L|no uncertainty reported|      5.00 keV       | Broad-band measurement|123615.19 +621009.0 (J2000)| Modelled datum|                                        |From reprocessed raw data; NED frequency assigned tomid-point of band in keV
2|0.5-8 keV (Chandra) | -15.80    ||log(erg/cm^2^/s)    |1.03E+18|  1.54E-11||Jy|2008ApJ...681.1163L|no uncertainty reported|      4.25 keV       | Broad-band measurement|123615.19 +621009.0 (J2000)| Modelled datum|                                        |From reprocessed raw data; NED frequency assigned tomid-point of band in keV
3|0.5-2 keV (Chandra) ||<-16.33    |log(erg/cm^2^/s)    |3.02E+17||1.55E-11|Jy|2008ApJ...681.1163L|no uncertainty reported|      1.25 keV       | Broad-band measurement|123615.19 +621009.0 (J2000)| Modelled datum|                                        |From reprocessed raw data; NED frequency assigned tomid-point of band in keV
4|B F435W (HST/ACS) AB      | 24.592    ||mag                 |6.98E+14|  5.29E-07||Jy|2007ApJ...660...81M|no uncertainty reported|    4297   A         | Broad-band measurement|12 36 15.208 +62 10 08.87 (J2000)| Flux integrated from map|                                        |From reprocessed raw data; Corrected for contaminatingsources
5|B (Subaru) AB       | 24.63     ||mag                 |6.77E+14|  5.11E-07||Jy|2006ApJ...653.1027W|no uncertainty reported| 4427.60   A         | Broad-band measurement|189.063367 62.169131 (J2000)| Flux in fixed aperture|3" diameter aperture                    |Averaged from previously published data
6|V (HST/ACS) AB      | 23.367    ||mag                 |5.08E+14|  1.63E-06||Jy|2007ApJ...660...81M|no uncertainty reported|    5907   A         | Broad-band measurement|12 36 15.208 +62 10 08.87 (J2000)| Flux integrated from map|                                        |From reprocessed raw data; Corrected for contaminatingsources
7|R (Keck II) AB      | 23.29     || mag                |4.62E+14|  1.75E-06||Jy|2004AJ....127.3121W|no uncertainty reported|   648.7   A         | Broad-band measurement|12 36 15.208 +62 10 08.87 (J2000)| Total flux|                                        |From new raw data
8|R (Subaru) AB       | 23.15     ||mag                 |4.59E+14|  1.99E-06||Jy|2006ApJ...653.1027W|no uncertainty reported| 6534.16   A         | Broad-band measurement|189.063367 62.169131 (J2000)| Flux in fixed aperture|3" diameter aperture                    |Averaged from previously published data
9|i F775W (HST/ACS) AB      | 22.090    ||mag                 |3.86E+14|  5.30E-06||Jy|2007ApJ...660...81M|no uncertainty reported|    7764   A         | Broad-band measurement|12 36 15.208 +62 10 08.87 (J2000)| Flux integrated from map|                                        |From reprocessed raw data; Corrected for contaminatingsources
10|I (Subaru) AB       | 22.20     ||mag                 |3.76E+14|  4.79E-06||Jy|2006ApJ...653.1027W|no uncertainty reported| 7975.89   A         | Broad-band measurement|189.063367 62.169131 (J2000)| Flux in fixed aperture|3" diameter aperture                    |Averaged from previously published data
11|z F850LP (HST/ACS) AB      | 21.425    ||mag                 |3.17E+14|  9.77E-06||Jy|2007ApJ...660...81M|no uncertainty reported|    9445   A         | Broad-band measurement|12 36 15.208 +62 10 08.87 (J2000)| Flux integrated from map|                                        |From reprocessed raw data; Corrected for contaminatingsources
12|HK' (QUIRC) AB      | 20.26     |+/-0.06 |mag                 |1.58E+14|  2.86E-05|+/-1.58E-06|Jy|2006ApJ...653.1027W|uncertainty|18947.38   A         | Broad-band measurement|189.063367 62.169131 (J2000)| Flux in fixed aperture|3" diameter aperture                    |Averaged from previously published data
13|3.6 microns (IRAC)  | 68.00     |+/-3.40 |microJy             |8.44E+13|  6.80E-05|+/-3.40E-06|Jy|2011AJ....141....1T|rms uncertainty|     3.550 microns   | Broad-band measurement|189.063309 62.169090 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
14|4.5 microns (IRAC)  | 52.20     |+/-2.61 |microJy             |6.67E+13|  5.22E-05|+/-2.61E-06|Jy|2011AJ....141....1T|rms uncertainty|     4.493 microns   | Broad-band measurement|189.063309 62.169090 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
15|5.8 microns (IRAC)  | 38.20     |+/-1.95 |microJy             |5.23E+13|  3.82E-05|+/-1.95E-06|Jy|2011AJ....141....1T|rms uncertainty|     5.731 microns   | Broad-band measurement|189.063309 62.169090 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
16|8.0 microns (IRAC)  | 46.10     |+/-2.36 |microJy             |3.81E+13|  4.61E-05|+/-2.36E-06|Jy|2011AJ....141....1T|rms uncertainty|     7.872 microns   | Broad-band measurement|189.063309 62.169090 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
17|16 microns (IRS)    | 311.0     |+/-12.2 |microJy             |1.90E+13|  3.11E-04|+/-1.22E-05|Jy|2011AJ....141....1T|rms uncertainty|      15.8 microns   | Broad-band measurement|189.063309 62.169090 (J2000)| From fitting to map|                                        |From new raw data
18|24 microns (MIPS)   | 325.9     |+/-5.3  |microJy             |1.27E+13|  3.26E-04|+/-5.30E-06|Jy|2011A&A...528A..35M|uncertainty|     23.68 microns   | Broad-band measurement|12 36 15.19 +62 10 08.66 (J2000)| Flux integrated from map|                                        |From new raw data
19|24 microns (MIPS)   | 325.0     |+/-6.6  |microJy             |1.27E+13|  3.25E-04|+/-6.60E-06|Jy|2011AJ....141....1T|rms uncertainty|     23.68 microns   | Broad-band measurement|189.063309 62.169090 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
1|MIPS 24 microns      | 327.      |+/-7.0  |microJy         |1.25E+13   |  327.E-06|+/-7.0E-06|Jy |1990IRASF.C...0000M|3sigma uncertainty| 25        microns   | Broad-band measurement|115813.1 +302058 (B1950)| Flux in fixed aperture|                                        |From new raw data
20|70 microns (MIPS)   | 4.9       |+/-0.3  |milliJy             |4.20E+12|  4.90E-03|+/-3.00E-04|Jy|2011A&A...528A..35M|uncertainty|     71.42 microns   | Broad-band measurement|12 36 15.19 +62 10 08.66 (J2000)| Flux integrated from map|                                        |From new raw data
2|70 microns (PACS)    | 4.5       |+/-0.6  |mJy             |4.283e+12  |  4.5E-03 |+/-0.6E-03|Jy |2.40e+01           |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
3|100 microns (PACS)   | 4.3       |+/-0.4  |mJy             |2.998e+12  |  4.3E-03 |+/-0.4E-03|Jy |2.40e+01           |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
4|160 microns (PACS)   | 9.2       |+/-1.0  |mJy             |1.874e+12  |  9.2E-03 |+/-1.0E-03|Jy |2.40e+01           |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
5|250 microns (SPIRE)  | 15.9      |+/-3.1  |mJy             |1.199e+12  |  15.9E-03|+/-3.1e-03|Jy |2.40e+01           |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
6|350 microns (SPIRE)  | 14.3      |+/-3.0  |mJy             |8.565e+11  |  14.3E-03|+/-3.0e-03|Jy |2.40e+01           |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
7|500 microns (SPIRE)  |           |<12.0   |mJy             |5.996e+11  |          |12.0e-03  |Jy |2.40e+01           |3sigma |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
8|1160 microns (Penner)|           |<1.7    |mJy             |2.58442E+11|          |1.7E-03   |Jy |2004MNRAS.354..779G|3sigma uncertainty|      1200 microns   | Broad-band measurement|16 36 55.9 +40 59 12 (J2000)| Flux integrated from map|S/N = 3.66                              |From new raw data
