
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-02-19T12:09:07PST



Photometric Data for SMM J140104.96+025223.5

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|2-8 keV (Chandra)   | |<5.8E-15   | erg/s/cm^2^        |1.21E+18| |4.79E-10|Jy|2008ApJ...675..262R|3 sigma|      5.00 keV       | Broad-band measurement|14 01 04.96 +02 52 24.8 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data; NED frequency assigned tomid-point of band in keV
2|0.5-8 keV (Chandra) | |<4.4E-15   | erg/s/cm^2^        |1.03E+18| |4.27E-10|Jy|2008ApJ...675..262R|3 sigma|      4.25 keV       | Broad-band measurement|14 01 04.96 +02 52 24.8 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data; NED frequency assigned tomid-point of band in keV
3|[O II] 3727         | 0.4E-16   |+/-0.1E-16|ergs cm^-2^ s^-1^   |8.04E+14|  4.98E-09|+/-1.24E-09|Jy|2006ApJ...651..713T|uncertainty|    3727   A         | Line measurement; flux integrated over line; lines measured in emission| | Flux integrated from map|From 2005AJ....129...53M                |Averaged from previously published data
4|H{beta}             | 0.3E-16   |+/-0.1E-16|ergs cm^-2^ s^-1^   |6.17E+14|  4.86E-09|+/-1.62E-09|Jy|2006ApJ...651..713T|uncertainty|    4861   A         | Line measurement; flux integrated over line; lines measured in emission| | Flux integrated from map|From 2005AJ....129...53M                |Averaged from previously published data
5|[O III] 4959        | |<0.2E-16   |ergs cm^-2^ s^-1^   |6.05E+14| |3.31E-09|Jy|2006ApJ...651..713T|no uncertainty reported|    4959   A         | Line measurement; flux integrated over line; lines measured in emission| | Flux integrated from map|From 2004ApJ...605L.109T                |Averaged from previously published data
6|[O III] 5007        | |<0.2E-16   |ergs cm^-2^ s^-1^   |5.99E+14| |3.34E-09|Jy|2006ApJ...651..713T|no uncertainty reported|    5007   A         | Line measurement; flux integrated over line; lines measured in emission| | Flux integrated from map|From 2005AJ....129...53M                |Averaged from previously published data
7|H{alpha} (IRTF)     | 1.2E-19   |+/-0.2E-19| W/m^2^             |4.57E+14|  2.63E-08|+/-4.38E-09|Jy|2004ApJ...617...64S|uncertainty|      6563 A         | Line measurement; flux integrated over line; lines measured in emission|140104.96 +025223.5 (J2000)| Flux integrated from map|                                        |From new raw data
8|H{alpha}            | 1.3E-16   |+/-0.4E-16|ergs cm^-2^ s^-1^   |4.57E+14|  2.84E-08|+/-8.75E-09|Jy|2006ApJ...651..713T|uncertainty|    6563   A         | Line measurement; flux integrated over line; lines measured in emission| | Flux integrated from map|From 2005AJ....129...53M                |Averaged from previously published data
9|3.6 microns (IRAC)  | 88        |+/-2    | microJy            |8.44E+13|  8.80E-05|+/-2.00E-06|Jy|2008ApJ...675..262R|uncertainty|     3.550 microns   | Broad-band measurement|14 01 04.96 +02 52 24.8 (J2000)| Flux in fixed aperture|                                        |From new raw data
10|4.5 microns (IRAC)  | 105       |+/-2    | microJy            |6.67E+13|  1.05E-04|+/-2.00E-06|Jy|2008ApJ...675..262R|uncertainty|     4.493 microns   | Broad-band measurement|14 01 04.96 +02 52 24.8 (J2000)| Flux in fixed aperture|                                        |From new raw data
11|5.6 microns (IRAC)  | 136       |+/-3    | microJy            |5.23E+13|  1.36E-04|+/-3.00E-06|Jy|2008ApJ...675..262R|uncertainty|     5.731 microns   | Broad-band measurement|14 01 04.96 +02 52 24.8 (J2000)| Flux in fixed aperture|                                        |From new raw data
12|8.0 microns (IRAC)  | 124       |+/-5    | microJy            |3.81E+13|  1.24E-04|+/-5.00E-06|Jy|2008ApJ...675..262R|uncertainty|     7.872 microns   | Broad-band measurement|14 01 04.96 +02 52 24.8 (J2000)| Flux in fixed aperture|                                        |From new raw data
13|24 microns (MIPS)   | 0.99      |+/-0.1  | milliJy            |1.27E+13|  9.90E-04|+/-1.00E-04|Jy|2008ApJ...675..262R|uncertainty|     23.68 microns   | Broad-band measurement|14 01 04.96 +02 52 24.8 (J2000)| From fitting to map|PSF fitting                             |From new raw data
13|24 microns (MIPS)   | 883.4     |+/-14.5  | uJy            |1.27E+13|  883.4E-06|+/-14.5E-06|Jy|2008ApJ...675..262R|uncertainty|     23.68 microns   | Broad-band measurement|14 01 04.96 +02 52 24.8 (J2000)| From fitting to map|PSF fitting                             |From new raw data
14|70 microns (MIPS)   | |<13        | milliJy            |4.20E+12| |1.30E-02|Jy|2008ApJ...675..262R|2sigma uncertainty reported|     71.42 microns   | Broad-band measurement|14 01 04.96 +02 52 24.8 (J2000)| Flux in fixed aperture|                                        |From new raw data
3|100 microns (PACS)   | 11.6      |+/-0.8  |mJy             |2.998e+12|11.6E-03|0.8E-03             |Jy|2005MNRAS.358..149P|3sigma uncertainty|     850   microns   | Broad-band measurement|12 37 11.7 +62 22 12 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
4|160 microns (PACS)  |  33.5      |+/-1.4 |mJy              |1.874e+12|33.5E-03|+/-1.4E-03  |Jy |2.40e+01          |3sigma|-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
5|250 microns (SPIRE)| 61.7      |+/-6.0 |mJy             |1.199e+12|61.7E-03|+/-6.0e-03 |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
15|350 microns (CSO)   | 75        |+/-10   |milliJy             |8.57E+11|  7.50E-02|+/-1.00E-02|Jy|2009ApJ...707..988W|rms noise|       350 microns   | Broad-band measurement|14 01 04.93 +02 52 24.1 (J2000)| Flux integrated from map|S/N=7.5 sigma                           |From new raw data
6|350 microns (SPIRE)| 63.1      |+/-3.8  |mJy             |8.565e+11|63.1E-03|+/-3.8e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
16|450 microns (SCUBA) | 6         |+/-8    |milliJy             |6.66E+11|  6.00E-03|+/-8.00E-03|Jy|2007MNRAS.376.1073Z|uncertainty|     450   microns   | Broad-band measurement|14 01 04.7 +02 52 28 (J2000)| Flux integrated from map|                                        |From reprocessed raw data
17|450 microns (SCUBA) | 42        |+/-7 |milliJy             |6.66E+11|  4.20E-02|+/-7.0E-03 |Jy|2002MNRAS.331..495S|no uncertainty reported|     450   microns   | Broad-band measurement|140105.0 +025225 (J2000)| Flux integrated from map|                                        |From new raw data
17|450 microns (SCUBA) | 41.9      |+/-6.9 |milliJy             |6.66E+11|  4.19E-02|+/-6.9E-03 |Jy|2002MNRAS.331..495S|no uncertainty reported|     450   microns   | Broad-band measurement|140105.0 +025225 (J2000)| Flux integrated from map|                                        |From new raw data
8|500 microns (SPIRE) | 48.5     |+/-4.0 |mJy             |5.996e+11|48.5E-03|+/-4.0e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
18|850 microns (SCUBA) | 13.4      |+/-1.4 |milliJy             |3.53E+11|  1.34E-02|+/-1.4E-03|Jy|2007MNRAS.376.1073Z|no uncertainty reported|     850   microns   | Broad-band measurement|14 01 04.7 +02 52 28 (J2000)| Flux integrated from map|S/N = 9.6                               |From reprocessed raw data
19|850 microns (SCUBA) | 12.3      |+/-1.7 |milliJy             |3.53E+11|  1.23E-02|+/-1.7E-03 |Jy|2002MNRAS.331..495S|no uncertainty reported|     850   microns   | Broad-band measurement|140105.0 +025225 (J2000)| Flux integrated from map|                                        |From new raw data
19|850 microns (SCUBA) | 14.6      |+/-1.8 |milliJy             |3.53E+11|  1.46E-02|+/-1.8E-03 |Jy|2002MNRAS.331..495S|no uncertainty reported|     850   microns   | Broad-band measurement|140105.0 +025225 (J2000)| Flux integrated from map|                                        |From new raw data
20|CO(1-0) (GBT)       | 0.4       |+/-0.05 |Jy km/s             |1.15E+11|  1.05E-07|+/-1.32E-08|Jy|2010ApJ...723.1139H|uncertainty|    115.27 GHz       | Line measurement; flux integrated over line; lines measured in emission|14 01 04.96 +02 52 23.5 (J2000)| Flux integrated from map|                                        |From new raw data
21|SCUBA 1350 microns  | 6.1       |+/-1.5 |milliJy             |2.22E+11|  6.1E-03|+/-1.5E-03|Jy|1999ApJ...519..610D|uncertainty| 1350      microns   | Broad-band measurement|164502.36 +462625.5 (J2000)| Flux integrated from map|                                        |From new raw data
14|1.4 GHz (VLA)       | 115.0     |+/-30.0| uJy                |1.40E+09|  115.0E-06|+/-30.0E-06|Jy|2004A&A...423..441B|uncertainty|    1.4    GHz       | Broad-band measurement|14 09 55.57 +56 28 26.47 (J2000)| Flux integrated from map|                                        |From new raw data
