
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-05-28T01:50:15PDT



Photometric Data for PJ105353.0, z=3.0053

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
4|UKIDSS J            | 0.24   |+/-0.001|mJy        |2.40161e+14|0.24E-3|+/-0.01E-3|Jy|2010Natur.464..733S|3rms uncertainty reported|      3344 A         | Broad-band measurement|21 35 11.6 -01 02 52.0 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
5|UKIDSS H            | 0.27   |+/-0.01|mJy         |1.83775e+14|0.27E-3|+/-0.01E-3|Jy|2010Natur.464..733S|3rms uncertainty reported|      3344 A         | Broad-band measurement|21 35 11.6 -01 02 52.0 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
6|UKIDSS K            | 0.22   |+/-0.01|mJy         |1.36207e+14|0.22E-3|+/-0.01E-3|Jy|2010Natur.464..733S|3rms uncertainty reported|      3344 A         | Broad-band measurement|21 35 11.6 -01 02 52.0 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
26|22 microns (WISE)  |        |<5.4|mJy            |1.36E+13||5.4E-03|Jy|2012AJ....144...49W|3sigma limit|        22 microns   | Broad-band measurement|213.942657 +11.495400 (J2000)| Not reported in paper|                                        |Averaged from previously published data
1|250 microns (SPIRE) | 1028.0     |+/-103.  |mJy         |1.199e+12|1028.0E-03 |+/-103.0e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
1|250 microns (SPIRE) | 1050.0     |+/-10.  |mJy         |1.199e+12|1050.0E-03 |+/-10.0e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
3|350 microns (SPIRE) | 996.0     |+/-100.  |mJy         |8.565e+11|996.0E-03 |+/-100.0e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
3|350 microns (SPIRE) | 1054.0     |+/-10.  |mJy         |8.565e+11|1054.0E-03 |+/-10.0e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
5|350 microns (PLANCK) | 2780.0    |+/-684.  |mJy        |8.57e+11|2780.0E-03 |+/-684.0e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
5|500 microns (SPIRE) | 735.0     |+/-74.  |mJy         |5.996e+11|735.0E-03 |+/-74.0e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
5|500 microns (SPIRE) | 777.0     |+/-7.  |mJy         |5.996e+11|777.0E-03 |+/-7.0e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
9|850 microns (SCUBA) | 198.0     |+/-11. |milliJy       |3.53E+11|  198.E-03|+/-11.E-03 |Jy|2002MNRAS.331..495S|no uncertainty reported|     850   microns   | Broad-band measurement|140105.0 +025225 (J2000)| Flux integrated from map|                                        |From new raw data
2|1.1mm (AzTEC)        | 98.0 |+/-10.| mJy  | 2.73E11| 98.0E-3| 10.0E-3 |Jy |2003MNRAS.343..293M|uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
5|GISMO(2000.0um)     |  19.0   |+/-2.0 |mJy          |150.000E+9|19.0E-03 |+/-2.0E-03|Jy|2010ApJ...709..210K|uncertainty|      870  microns   | Broad-band measurement|16 35 55.67 +66 12 59.51 (J2000)| Flux integrated from map|                                        |From new raw data
21|1.4GHz (VLA)       |   6.5 |+/-1.3|mJy| 1.4E9   |6.5E-03 |1.3E-03 |Jy |2003MNRAS.343..293M|3rms uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
21|1.4GHz (VLA)       |   2.26 |+/-0.14|mJy| 1.4E9   |2.26E-03 |0.14E-03 |Jy |2003MNRAS.343..293M|3rms uncertainty|    4.25   keV       | Broad-band measurement|16 36 55.79 +40 59 10.5 (J2000)| Flux integrated from map|                                        |From new raw data; NED frequency assigned to mid-point ofband in keV
