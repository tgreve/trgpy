
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-04-03T14:24:27PDT



Photometric Data for ABELL 2218 ARC L

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|2-8 keV (Chandra)   | |<2.8E-15   | erg/s/cm^2^        |1.21E+18| |2.31E-10|Jy|2008ApJ...675..262R|3 sigma|      5.00 keV       | Broad-band measurement|16 35 55.16 +66 11 50.8 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data; NED frequency assigned tomid-point of band in keV
2|0.5-8 keV (Chandra) | |<2.1E-15   | erg/s/cm^2^        |1.03E+18| |2.04E-10|Jy|2008ApJ...675..262R|3 sigma|      4.25 keV       | Broad-band measurement|16 35 55.16 +66 11 50.8 (J2000)| Flux in fixed aperture|                                        |From reprocessed raw data; NED frequency assigned tomid-point of band in keV
3|F606W (HST/WFPC2)   | 20.25     |+/-0.02 |mag                 |5.05E+14|  2.70E-05|+/-4.98E-07|Jy|2005ApJ...627...32S|uncertainty|    5934   A         | Broad-band measurement| | Flux integrated from map|                                        |From new raw data
4|3.5 microns (IRAC)  | 182       |+/-4    | microJy            |8.44E+13|  1.82E-04|+/-4.00E-06|Jy|2008ApJ...675..262R|uncertainty|     3.550 microns   | Broad-band measurement|16 35 55.16 +66 11 50.8 (J2000)| Flux in fixed aperture|                                        |From new raw data
5|4.5 microns (IRAC)  | 147       |+/-3    | microJy            |6.67E+13|  1.47E-04|+/-3.00E-06|Jy|2008ApJ...675..262R|uncertainty|     4.493 microns   | Broad-band measurement|16 35 55.16 +66 11 50.8 (J2000)| Flux in fixed aperture|                                        |From new raw data
6|5.7 microns (IRAC)  | 107       |+/-3    | microJy            |5.23E+13|  1.07E-04|+/-3.00E-06|Jy|2008ApJ...675..262R|uncertainty|     5.731 microns   | Broad-band measurement|16 35 55.16 +66 11 50.8 (J2000)| Flux in fixed aperture|                                        |From new raw data
7|8.0 microns (IRAC)  | 107       |+/-5    | microJy            |3.81E+13|  1.07E-04|+/-5.00E-06|Jy|2008ApJ...675..262R|uncertainty|     7.872 microns   | Broad-band measurement|16 35 55.16 +66 11 50.8 (J2000)| Flux in fixed aperture|                                        |From new raw data
8|24 microns (MIPS)   | 1.67      |+/-0.1  | milliJy            |1.27E+13|  1.67E-03|+/-1.00E-04|Jy|2008ApJ...675..262R|uncertainty|     23.68 microns   | Broad-band measurement|16 35 55.16 +66 11 50.8 (J2000)| From fitting to map|PSF fitting                             |From new raw data
9|70 microns (MIPS)   | 7.4       |+/-1.5  | milliJy            |4.20E+12|  7.40E-03|+/-1.50E-03|Jy|2008ApJ...675..262R|uncertainty|     71.42 microns   | Broad-band measurement|16 35 55.16 +66 11 50.8 (J2000)| Flux in fixed aperture|                                        |From new raw data
10|450 microns (SCUBA) | 17.1      |+/-5.1  | milliJy            |6.66E+11|  1.71E-02|+/-5.10E-03|Jy|2008MNRAS.384.1611K|rms uncertainty|       450 microns   | Broad-band measurement|163555.2 +661150 (J2000)| Flux integrated from map|S/N = 4.7                               |From new raw data
11|450 microns (SCUBA) | 29.1      |+/-8.7  |milliJy             |6.66E+11|  2.91E-02|+/-8.70E-03|Jy|2006MNRAS.368..487K|uncertainty|     450   microns   | Broad-band measurement|163555.2 +661150 (J2000)| Flux integrated from map|                                        |From new raw data
12|850 microns (SCUBA) | 3.1       |+/-0.7  | milliJy            |3.53E+11|  3.10E-03|+/-7.00E-04|Jy|2008MNRAS.384.1611K|rms uncertainty|       850 microns   | Broad-band measurement|163555.2 +661150 (J2000)| Flux integrated from map|S/N = 3.8                               |From new raw data
13|850 microns (SCUBA) | 3.1       |+/-0.7  |milliJy             |3.53E+11|  3.10E-03|+/-7.00E-04|Jy|2006MNRAS.368..487K|uncertainty|     850   microns   | Broad-band measurement|163555.2 +661150 (J2000)| Flux integrated from map|                                        |From new raw data
14|CO(2-1) (IRAM)      | 1.2       |+/-0.2  | Jy km/s            |2.31E+11|  9.68E-07|+/-1.61E-07|Jy|2009A&A...496...45K|uncertainty|   230.538 GHz       | Line measurement; flux integrated over line; lines measured in emission|16 35 55.05 +66 11 50.7 (J2000)| Flux integrated from map|                                        |From new raw data
15|3 mm (IRAM)         | |<1.4       | milliJy            |9.99E+10| |1.40E-03|Jy|2009A&A...496...45K|3sigma uncertainty|         3 mm        | Broad-band measurement|16 35 55.05 +66 11 50.7 (J2000)| Flux integrated from map|                                        |From new raw data
