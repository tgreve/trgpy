
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-06-16T17:14:05PDT



Photometric Data for [HB89] 2343+125:BX0442

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|G (WHT)             | 24.48     ||mag                 |6.38E+14|  5.86E-07||Jy|2006ApJ...647..128E|no uncertainty reported|    0.47   microns   | Broad-band measurement|| Flux in fixed aperture|                                        |Averaged from previously published data
2|H{alpha} (Keck II)  | 7.1E-17   |+/-0.3E-17|erg s^-1^ cm^-2^    |4.57E+14|  7.10E+06|+/-3.00E+05|Jy-Hz|2006ApJ...646..107E|uncertainty|    6563   A         | Line measurement; flux integrated over line; lines measured in emission|23 46 19.36 +12 47 59.69 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
3|J (Hale/WIRC)       | 22.21     ||mag                 |2.40E+14|  2.04E-06||Jy|2006ApJ...646..107E|no uncertainty reported|    1.25   microns   | Broad-band measurement|23 46 19.36 +12 47 59.69 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data; derived from aflux in a different band and a color
4|K_s (Hale/WIRC)     | 19.85     ||mag                 |1.39E+14|  7.69E-06||Jy|2006ApJ...646..107E|no uncertainty reported|    2.15   microns   | Broad-band measurement|23 46 19.36 +12 47 59.69 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data
5|CO(3-2) (PdBI)      ||<0.08      |Jy km/s             |3.46E+11|  1.56E+05|2.90E+04|Jy-Hz|2010Natur.463..781T|3 sigma|   345.998 GHz       | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|                                        |From new raw data
