
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-06-17T09:40:16PDT



Photometric Data for SDF J132415.7+273058

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
11|CARMA 165GHz      |      |<0.17 |mJy                 |1.65E+11|  |0.17E-03|Jy|2011ApJ...736L..28C|1sigma uncertainty|     13006 A         | Broad-band measurement|| Flux in fixed aperture|                                        |From new raw data
