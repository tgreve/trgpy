
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-07-10T13:42:15PDT



Photometric Data for SPT-SJ214654-5507.8

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
5|250 microns (SPIRE)| 43.      |+/-10.0 |mJy             |1.199e+12| 43.0E-03|+/-10.0e-03 |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
6|350 microns (SPIRE)| 72.      |+/-11.  |mJy             |8.565e+11|72.E-03 |+/-11.0e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
8|500 microns (SPIRE) | 108.     |+/-15. |mJy             |5.996e+11|108.0E-03 |+/-15.0e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
1|870 microns (LABOCA)| 70.0     |+/-13.  |milliJy        |3.45E+11|  70.0E-03|+/-13.0E-03|Jy|2009ApJ...707.1201W|uncertainty|       870 microns   | Broad-band measurement|03 32 29.33 -27 56 19.3 (J2000)| Flux integrated from map|S/N = 4.6                               |From new raw data
1|1.4 mm (SPT)        | 28.5     |+/-8.1 |milliJy         |2.20E+11|  28.5E-03|+/-8.1E-03|Jy|2010ApJ...719..763V|uncertainty|       1.4 mm        | Broad-band measurement|74.804 -59.708 (J2000)| Flux integrated from map|De-boosted flux; S/N = 7.05             |From new raw data
3|2.0 mm (SPT)        | 8.1     |+/-1.4 |milliJy          |1.50E+11|  8.1E-03|+/-1.4E-03|Jy|2010ApJ...719..763V|uncertainty|       2.0 mm        | Broad-band measurement|74.804 -59.708 (J2000)| Flux integrated from map|De-boosted flux; S/N = 6.20             |From new raw data
1|3.0mm (ALMA)        | 0.99 | 0.16 |milliJy            |1.0E+11| 0.99E-3 |0.16E-3 |Jy|2007MNRAS.376.1073Z|no uncertainty reported|     850   microns   | Broad-band measurement|02 39 51.9 -01 35 55 (J2000)| Flux integrated from map|S/N = 19.9                              |From reprocessed raw data
3|41.9GHz (ATCA)      |         |<135.0|microJy             |41.9E+09||135.0E-06|Jy|2010ApJ...719..763V|3sigma uncertainty|       2.0 mm        | Broad-band measurement|74.804 -59.708 (J2000)| Flux integrated from map|De-boosted flux; S/N = 6.20             |From new raw data
