
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-05-03T03:12:46PDT



Photometric Data for SMM J023951.87-013558.8

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|3.6 microns (IRAC)  | 9.8290E+01|+/-8.5146E-02|microJy             |8.44E+13|  9.83E-05|+/-8.51E-08|Jy|2013SSTSLC4.2....0C|uncertainty|3.55       microns   | Broad-band measurement|| Flux in fixed aperture|5.8" aperture                           |From new raw data
2|3.6 microns (IRAC)  | 7.7237E+01|+/-6.9348E-02|microJy             |8.44E+13|  7.72E-05|+/-6.93E-08|Jy|2013SSTSLC4.2....0C|uncertainty|3.55       microns   | Broad-band measurement|| Flux in fixed aperture|3.8" aperture                           |From new raw data
3|4.5 microns (IRAC)  | 1.1107E+02|+/-8.9364E-02|microJy             |6.67E+13|  1.11E-04|+/-8.94E-08|Jy|2013SSTSLC4.2....0C|uncertainty|4.493      microns   | Broad-band measurement|| Flux in fixed aperture|3.8" aperture                           |From new raw data
4|4.5 microns (IRAC)  | 1.3815E+02|+/-1.2532E-01|microJy             |6.67E+13|  1.38E-04|+/-1.25E-07|Jy|2013SSTSLC4.2....0C|uncertainty|4.493      microns   | Broad-band measurement|| Flux in fixed aperture|5.8" aperture                           |From new raw data
5|5.8 microns (IRAC)  | 1.9915E+02|+/-4.6486E-01|microJy             |5.23E+13|  1.99E-04|+/-4.65E-07|Jy|2013SSTSLC4.2....0C|uncertainty|5.731      microns   | Broad-band measurement|| Flux in fixed aperture|5.8" aperture                           |From new raw data
6|5.8 microns (IRAC)  | 1.7725E+02|+/-3.4786E-01|microJy             |5.23E+13|  1.77E-04|+/-3.48E-07|Jy|2013SSTSLC4.2....0C|uncertainty|5.731      microns   | Broad-band measurement|| Flux in fixed aperture|3.8" aperture                           |From new raw data
3|IRAS 12 microns     | |<91        |milliJy             |2.50E+13| |91.0E-03|Jy|1999ApJ...519..610D|3sisgma uncertainty reported| 12        microns   | Broad-band measurement|164502.36 +462625.5 (J2000)| Integrated from scans|                                        |Averaged from previously published data
4|ISOCAM 15 microns  | 1.2    |+/-0.4  |milliJy             |2.07E+13|  1.2E-03|+/-0.4E-03|Jy|1997MNRAS.289..465G|estimated error|14.5       microns   | Broad-band measurement|123634.37 +621238.6 (J2000)| Flux integrated from map|                                        |From new raw data
5|24 microns (MIPS)   | 1.24      |+/-10  %|milliJy             |1.27E+13|  1.24E-03|+/-1.24E-04 |Jy|2009A&A...502..541E|uncertainty|     23.68 microns   | Broad-band measurement| | Flux in fixed aperture|                                        |From reprocessed raw data
6|IRAS 25 microns     | |<85        |milliJy             |1.20E+13| |85.0E-03|Jy|1999ApJ...519..610D|3sisgma uncertainty reported| 25        microns   | Broad-band measurement|164502.36 +462625.5 (J2000)| Integrated from scans|                                        |Averaged from previously published data
2|29.3microns (monochromatic)   | 1.44      |+/-0.3 |milliJy             |1.02E+13|  1.44E-03|+/-0.3E-03 |Jy|2007ApJ...660.1060V|1sigma uncertainty reported|     7.7   microns   | Broad-band measurement|02 39 51.87 -01 35 58.8 (J2000)| Flux integrated from map|                                        |From new raw data
7|IRAS 60 microns     | |<428        |milliJy             |5.00E+12| |428.0E-03|Jy|1999ApJ...519..610D|3sisgma uncertainty reported| 60        microns   | Broad-band measurement|164502.36 +462625.5 (J2000)| Integrated from scans|                                        |Averaged from previously published data
9|70 microns (MIPS)   | 15        |+/-30  % |milliJy             |4.20E+12|  1.50E-02|+/-4.5E-03 |Jy|2009A&A...502..541E|uncertainty reported|     71.42 microns   | Broad-band measurement| | Flux in fixed aperture|Tentative detection                     |From reprocessed raw data
8|IRAS 100 microns    | |<715       |milliJy             |3.00E+12| |715.0E-03|Jy|1999ApJ...519..610D|3sisgma uncertainty reported| 100       microns   | Broad-band measurement|164502.36 +462625.5 (J2000)| Integrated from scans|                                        |Averaged from previously published data
10|160 microns (MIPS)  | 16        |+/-30  % |milliJy             |1.92E+12|  1.60E-02|+/-4.8E-03 |Jy|2009A&A...502..541E|uncertainty reported|     155.9 microns   | Broad-band measurement| | Flux in fixed aperture|                                        |From reprocessed raw data
11|350 microns (CSO/SHARC-II)   | 29        |+/-9    |milliJy             |8.57E+11|  2.90E-02|+/-9.00E-03|Jy|2009ApJ...707..988W|1sigma noise|       350 microns   | Broad-band measurement|02 39 51.90 -01 35 58.8 (J2000)| Flux integrated from map|S/N=3.1 sigma                           |From new raw data
12|350 microns (SCUBA) |           |<323.0  |milliJy             |8.573E+11| |323.0E-03|Jy|2007MNRAS.376.1073Z|3sigma uncertainty|     450   microns   | Broad-band measurement|02 39 51.9 -01 35 55 (J2000)| Flux integrated from map|                                        |From reprocessed raw data
13|450 microns (SCUBA) | -2        |+/-19   |milliJy             |6.66E+11| -2.00E-03|+/-1.90E-02|Jy|2007MNRAS.376.1073Z|1sigma uncertainty|     450   microns   | Broad-band measurement|02 39 51.9 -01 35 55 (J2000)| Flux integrated from map|                                        |From reprocessed raw data
14|450 microns (SCUBA) | 85        |+/-10 |milliJy             |6.66E+11|  8.50E-02|+/-10.E-03 |Jy|2002MNRAS.331..495S|no uncertainty reported|     450   microns   | Broad-band measurement|023951.9 -013559 (J2000)| Flux integrated from map|                                        |From new raw data
15|450 microns (SCUBA) | 69        |+/-15 |milliJy             |6.66E+11|  6.90E-02|+/-15.E-03 |Jy|2002MNRAS.331..495S|no uncertainty reported|     450   microns   | Broad-band measurement|023951.9 -013559 (J2000)| Flux integrated from map|                                        |From new raw data
16|750 microns (SCUBA) | 28.0      |+/-5.0 |milliJy             |3.99E+11|  28.0E-03|+/-5.0E-03 |Jy|2007MNRAS.376.1073Z|no uncertainty reported|     850   microns   | Broad-band measurement|02 39 51.9 -01 35 55 (J2000)| Flux integrated from map|S/N = 19.9                              |From reprocessed raw data
17|850 microns (SCUBA) | 20.5      |+/-1.9 |milliJy             |3.53E+11|  2.05E-02|+/-1.9E-03 |Jy|2002MNRAS.331..495S|no uncertainty reported|     850   microns   | Broad-band measurement|023951.9 -013559 (J2000)| Flux integrated from map|                                        |From new raw data
18|850 microns (SCUBA) | 23.0      |+/-1.9 |milliJy             |3.53E+11|  2.30E-02|+/-1.9E-03 |Jy|2002MNRAS.331..495S|no uncertainty reported|     850   microns   | Broad-band measurement|023951.9 -013559 (J2000)| Flux integrated from map|                                        |From new raw data
19|850 microns (SCUBA) | 26.0      |+/-3.0 |milliJy             |3.53E+11|  2.60E-02|+/-3.0E-03 |Jy|2002MNRAS.331..495S|no uncertainty reported|     850   microns   | Broad-band measurement|023951.9 -013559 (J2000)| Flux integrated from map|                                        |From new raw data
20|1270 microns (PDBI) | 7.0      |+/-1.2 |milliJy             |2.35E+11|  7.0E-03|+/-1.2E-03 |Jy|2002MNRAS.331..495S|no uncertainty reported|     850   microns   | Broad-band measurement|023951.9 -013559 (J2000)| Flux integrated from map|                                        |From new raw data
21|SCUBA 1350 microns  | 5.7      |+/-1.0 |milliJy             |2.22E+11|  5.7E-03|+/-1.0E-03|Jy|1999ApJ...519..610D|uncertainty| 1350      microns   | Broad-band measurement|164502.36 +462625.5 (J2000)| Flux integrated from map|                                        |From new raw data
22|212.537 GHz (PdBI)  | 6.2       |+/-0.2  |milliJy             |2.13E+11|  6.20E-03|+/-2.00E-04|Jy|2011ApJ...730...18W|uncertainty|   212.537 GHz       | Broad-band measurement|02 38 51.87 -01 35 58.8 (J2000)| Flux integrated from map|Flux includes the CI(2-1) line          |From new raw data
23|SCUBA 2000 microns  |      |<8.4 |milliJy             |1.49896e+11| |8.4E-03|Jy|1999ApJ...519..610D|3rms uncertainty| 1350      microns   | Broad-band measurement|164502.36 +462625.5 (J2000)| Flux integrated from map|                                        |From new raw data
24|129.244 GHz (PdBI)  | |<0.5       |milliJy             |1.29E+11| |5.00E-04|Jy|2011ApJ...730...18W|3sigma|   129.244 GHz       | Broad-band measurement|02 38 51.87 -01 35 58.8 (J2000)| Flux integrated from map|                                        |From new raw data
25|32.3 GHz (EVLA)     | |<60.  | microJy            |32.3E+09| |60.E-06|Jy|2007MNRAS.380..199I|2 rms uncertainty|       1.4 GHz       | Broad-band measurement|10 52 28.995 +57 22 22.42 (J2000)| Flux integrated from map|                                        |From reprocessed raw data
26|32.0 GHz (JVLA)     |57.0       |+/-25.  | microJy            |32.0E+09|57.0E-06|+/-25.E-06|Jy|2007MNRAS.380..199I|2 rms uncertainty|       1.4 GHz       | Broad-band measurement|10 52 28.995 +57 22 22.42 (J2000)| Flux integrated from map|                                        |From reprocessed raw data
27|8.7 GHz (VLA)       |       |<57.0  | microJy            |8.7E+09|  |57.0E-06|Jy|2007MNRAS.380..199I|3 rms uncertainty|       1.4 GHz       | Broad-band measurement|10 52 28.995 +57 22 22.42 (J2000)| Flux integrated from map|                                        |From reprocessed raw data
28|5.0 GHz (VLA)       | 130.      |+/-22.  | microJy            |5.00E+09|  130.E-06|+/-22.E-06|Jy|2007MNRAS.380..199I|rms uncertainty|       1.4 GHz       | Broad-band measurement|10 52 28.995 +57 22 22.42 (J2000)| Flux integrated from map|                                        |From reprocessed raw data
29|1.4 GHz (VLA)       | 526.      |+/-10.  | microJy            |1.40E+09|  526.E-06|+/-10.E-06|Jy|2007MNRAS.380..199I|rms uncertainty|       1.4 GHz       | Broad-band measurement|10 52 28.995 +57 22 22.42 (J2000)| Flux integrated from map|                                        |From reprocessed raw data
