
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-05-28T01:42:09PDT



Photometric Data for SPT-S233227-5358.5, z=2.738

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|352 microns (APEX) | 425       |+/-39   |mJy             |8.52E+11|  425.0E-03|+/-39.0E-03|Jy|2010Natur.464..733S|uncertainty|       352 microns   | Broad-band measurement|21 35 11.6 -01 02 52.0 (J2000)| Flux in fixed aperture|                                        |From new raw data
2|870 microns (APEX) | 150       |+/-11   |mJy             |3.45E+11|  150.0E-03|+/-11.0E-03|Jy|2010Natur.464..733S|uncertainty|       870 microns   | Broad-band measurement|21 35 11.6 -01 02 52.0 (J2000)| Flux in fixed aperture|                                        |From new raw data
3|1360 microns (SPT) | 34.4      | 4.7    |mJy             |2.20436E+11| 34.4E-3 |4.7E-3 |Jy|2007MNRAS.376.1073Z|no uncertainty reported|     850   microns   | Broad-band measurement|02 39 51.9 -01 35 55 (J2000)| Flux integrated from map|S/N = 19.9                              |From reprocessed raw data
4|0.85cm (VLA)       |           |<120|microJy             |35.0E+09| |120.0E-06|Jy|2010A&A...518L..35I|3rms uncertainty|      4.49 cm        | Broad-band measurement| | Flux integrated from map|                                        |From new raw data
5|0.97cm (VLA)       |           |<120|microJy             |31.0E+09| |120.0E-06|Jy|2010A&A...518L..35I|3rms uncertainty|      4.49 cm        | Broad-band measurement| | Flux integrated from map|                                        |From new raw data
