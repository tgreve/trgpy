\queryDateTime = 2018-11-27T11:31:53PST
\source = /hydra/workarea/irsaviewer/temp_files/IpacTableFromSource3921649364618972268.tbl
\QUERY_STATUS = OK
\CatalogTargetColName = Coordinates Targeted
\Description = Published and Homogenized [Frequency, Flux Dens...
\LINK = http://ned.ipac.caltech.edu/cgi-bin/datasearch?sea
\
z=0.01594
|No.   |Observed Passband   |Photometry Measurement|Uncertainty  |Units               |Frequency|Flux Density|Upper limit of uncertainty|Lower limit of uncertainty|Upper limit of Flux Density|Lower limit of Flux Density|NED Uncertainty|NED Units|Refcode            |Significance           |Published frequency|Frequency Mode                                                         |Coordinates Targeted            |Spatial Mode                                            |Qualifiers                             |Comments                                                                                                                                                           |
|int   |char                |double                |char         |char                |double   |double      |double                    |double                    |double                     |double                     |char           |char     |char               |char                   |char               |char                                                                   |char                            |char                                                    |char                                   |char                                                                                                                                                               |
|      |                    |                      |             |                    |Hz       |Jy          |                          |                          |                           |                           |               |         |                   |                       |                   |                                                                       |                                |                                                        |                                       |                                                                                                                                                                   |
|      |                    |                      |             |                    |         |            |                          |                          |                           |                           |               |         |                   |                       |                   |                                                                       |                                |                                                        |                                       |                                                                                                                                                                   |
 1     |2-10 keV (ASCA)     |3.6E-13               |             |ergs/s/cm^2^        |1.45E+18 |2.48E-08    |                          |                          |                           |                           |               |Jy       |2001ApJS..133....1U|no uncertainty reported|6.00 keV           |Broad-band measurement                                                 |068.5087 -08.5895 (J2000)       |Flux integrated from map                                |                                       |From reprocessed raw data; Extinction-corrected for MilkyWay; NED frequency assigned to mid-point of band in keV                                                   
 2     |2-10 keV (XMM)      |2.8E-13               |+/-4.2E-14   |erg/cm^2^/s         |1.45E+18 |1.90E-08    |2.9E-09                   |2.9E-09                   |                           |                           |+/-2.90E-09    |Jy       |2011A&A...535A..93P|uncertainty            |6.00 keV           |Broad-band measurement                                                 |                                |Modelled datum                                          |                                       |From new raw data; NED frequency assigned to mid-point ofband in keV                                                                                               
 3     |2-10 keV (XMM)      |2.6E-13               |             |erg/s/cm^2^         |1.45E+18 |1.79E-08    |                          |                          |                           |                           |               |Jy       |2011MNRAS.413.1206B|no uncertainty reported|6.00 keV           |Broad-band measurement                                                 |068.501 -08.579 (J2000)         |Modelled datum                                          |                                       |From reprocessed raw data; NED frequency assigned tomid-point of band in keV                                                                                       
 4     |0.7-7 keV (ASCA)    |4.8E-13               |             |ergs/s/cm^2^        |9.31E+17 |5.16E-08    |                          |                          |                           |                           |               |Jy       |2001ApJS..133....1U|no uncertainty reported|3.85 keV           |Broad-band measurement                                                 |068.5087 -08.5895 (J2000)       |Flux integrated from map                                |                                       |From reprocessed raw data; Extinction-corrected for MilkyWay; NED frequency assigned to mid-point of band in keV                                                   
 5     |0.2-4 keV (EINSTEIN)|6.5E-13               |             |ergs sec^-1^ cm^-2^ |5.25E+17 |1.24E-07    |                          |                          |                           |                           |               |Jy       |1992ApJS...80..531F|no uncertainty reported|2.1    keV         |Broad-band measurement; synthetic band                                 |04 31 35 -08 40 53 (B1950)      |Flux integrated from map                                |                                       |From reprocessed raw data; Extinction-corrected for MilkyWay; NED frequency assigned to mid-point of band in keV                                                   
 6     |0.7-2 keV (ASCA)    |2.0E-13               |             |ergs/s/cm^2^        |3.26E+17 |6.13E-08    |                          |                          |                           |                           |               |Jy       |2001ApJS..133....1U|no uncertainty reported|1.35 keV           |Broad-band measurement                                                 |068.5087 -08.5895 (J2000)       |Flux integrated from map                                |                                       |From reprocessed raw data; Extinction-corrected for MilkyWay; NED frequency assigned to mid-point of band in keV                                                   
 7     |0.5-2 keV (XMM)     |1.8E-13               |+/-2.4E-14   |erg/cm^2^/s         |3.02E+17 |5.86E-08    |8.0E-09                   |8.0E-09                   |                           |                           |+/-7.95E-09    |Jy       |2011A&A...535A..93P|uncertainty            |1.25 keV           |Broad-band measurement                                                 |                                |Modelled datum                                          |                                       |From new raw data; NED frequency assigned to mid-point ofband in keV                                                                                               
 8     |1482A (IUE)         |5.6E-15               |+/-0.22E-14  |ergs cm^-2 s^-1 A^-1|2.02E+15 |4.11E-04    |1.6E-04                   |1.6E-04                   |                           |                           |+/-1.61E-04    |Jy       |1993ApJS...86....5K|uncertainty            |1482   A           |Broad-band measurement; flux integrated over line                      |                                |Flux in fixed aperture                                  |20"x10" aperture                       |Averaged from new and transformed previously published data                                                                                                        
 9     |1913A (IUE)         |4.3E-15               |+/-0.08E-14  |ergs cm^-2 s^-1 A^-1|1.57E+15 |5.26E-04    |9.8E-05                   |9.8E-05                   |                           |                           |+/-9.78E-05    |Jy       |1993ApJS...86....5K|uncertainty            |1913   A           |Broad-band measurement; flux integrated over line                      |                                |Flux in fixed aperture                                  |20"x10" aperture                       |Averaged from new and transformed previously published data                                                                                                        
 10    |UVW2 (Swift) AB     |1.5E+01               |+/-0.10      |mag                 |1.48E+15 |5.19E-03    |4.8E-04                   |4.8E-04                   |                           |                           |+/-4.78E-04    |Jy       |2014ApJS..212...18B|uncertainty            |2026   A           |Broad-band measurement                                                 |68.50016000 -8.57923000 (J2000) |Flux in fixed aperture                                  |80"x60" aperture                       |From new raw data; Extinction-corrected for Milky Way                                                                                                              
 11    |UVW2 (Swift) AB     |1.6E+01               |+/-0.10      |mag                 |1.48E+15 |1.60E-03    |1.5E-04                   |1.5E-04                   |                           |                           |+/-1.48E-04    |Jy       |2014ApJS..212...18B|uncertainty            |2026   A           |Broad-band measurement                                                 |68.50016000 -8.57923000 (J2000) |Flux in fixed aperture                                  |80"x60" aperture                       |From new raw data                                                                                                                                                  
 12    |UVW2 (XMM-OM)       |9.3E-01               |             |milliJy             |1.41E+15 |9.30E-04    |                          |                          |                           |                           |               |Jy       |2011A&A...535A..93P|no uncertainty reported|2120 A             |Broad-band measurement                                                 |                                |Flux in fixed aperture                                  |                                       |From new raw data                                                                                                                                                  
 13    |UVM2 (Swift) AB     |1.5E+01               |+/-0.10      |mag                 |1.34E+15 |4.92E-03    |4.5E-04                   |4.5E-04                   |                           |                           |+/-4.53E-04    |Jy       |2014ApJS..212...18B|uncertainty            |2239   A           |Broad-band measurement                                                 |68.50016000 -8.57923000 (J2000) |Flux in fixed aperture                                  |80"x60" aperture                       |From new raw data; Extinction-corrected for Milky Way                                                                                                              
 14    |UVM2 (Swift) AB     |1.6E+01               |+/-0.10      |mag                 |1.34E+15 |1.45E-03    |1.3E-04                   |1.3E-04                   |                           |                           |+/-1.34E-04    |Jy       |2014ApJS..212...18B|uncertainty            |2239   A           |Broad-band measurement                                                 |68.50016000 -8.57923000 (J2000) |Flux in fixed aperture                                  |80"x60" aperture                       |From new raw data                                                                                                                                                  
 15    |UVW1 (Swift) AB     |1.5E+01               |+/-0.10      |mag                 |1.15E+15 |2.38E-03    |2.2E-04                   |2.2E-04                   |                           |                           |+/-2.19E-04    |Jy       |2014ApJS..212...18B|uncertainty            |2598   A           |Broad-band measurement                                                 |68.50016000 -8.57923000 (J2000) |Flux in fixed aperture                                  |80"x60" aperture                       |From new raw data                                                                                                                                                  
 16    |UVW1 (Swift) AB     |1.5E+01               |+/-0.10      |mag                 |1.15E+15 |5.69E-03    |5.2E-04                   |5.2E-04                   |                           |                           |+/-5.24E-04    |Jy       |2014ApJS..212...18B|uncertainty            |2598   A           |Broad-band measurement                                                 |68.50016000 -8.57923000 (J2000) |Flux in fixed aperture                                  |80"x60" aperture                       |From new raw data; Extinction-corrected for Milky Way                                                                                                              
 17    |u (SDSS) AB         |1.4E+01               |+/-0.05      |mag                 |8.44E+14 |1.10E-02    |5.1E-04                   |5.1E-04                   |                           |                           |+/-5.07E-04    |Jy       |2014ApJS..212...18B|uncertainty            |3551   A           |Broad-band measurement                                                 |68.50016000 -8.57923000 (J2000) |Flux in fixed aperture                                  |80"x60" aperture                       |From new raw data; Extinction-corrected for Milky Way                                                                                                              
 18    |u (SDSS) AB         |1.5E+01               |+/-0.05      |mag                 |8.44E+14 |5.76E-03    |2.7E-04                   |2.7E-04                   |                           |                           |+/-2.65E-04    |Jy       |2014ApJS..212...18B|uncertainty            |3551   A           |Broad-band measurement                                                 |68.50016000 -8.57923000 (J2000) |Flux in fixed aperture                                  |80"x60" aperture                       |From new raw data                                                                                                                                                  
 19    |U_T (VATT)          |1.4E+01               |+/-0.014     |mag                 |8.19E+14 |7.15E-03    |9.5E-05                   |9.5E-05                   |                           |                           |+/-9.49E-05    |Jy       |2005ApJ...630..784T|uncertainty            |3660   A           |Broad-band measurement                                                 |04 33 59.20 -08 35 56.3 (J2000) |Total flux                                              |                                       |From new raw data; derived from a flux in a different bandand a color; Standard Johnson UBVRI filters assumed                                                      
 20    |U (U_T)             |1.4E+01               |+/-0.13      |mag                 |8.19E+14 |6.45E-03    |8.4E-04                   |8.4E-04                   |                           |                           |+/-8.44E-04    |Jy       |1991RC3.9.C...0000d|rms uncertainty        |3660       A       |Broad-band measurement                                                 |043135.5 -084042 (B1950)        |From multi-aperture data                                |                                       |Homogenized from new and previously published data; StandardJohnson UBVRI filters assumed                                                                          
 21    |U (U_T^0)           |1.3E+01               |             |mag                 |8.19E+14 |9.50E-03    |                          |                          |                           |                           |               |Jy       |1991RC3.9.C...0000d|no uncertainty reported|3660       A       |Broad-band measurement                                                 |043135.5 -084042 (B1950)        |From multi-aperture data                                |                                       |Homogenized from new and previously published data;Extinction-corrected for internal and Milky Way and K-correction applied; Standard Johnson UBVRI filters assumed
 23    |103a-O (POSS-I O)   |1.6E+01               |             |mag                 |7.40E+14 |1.01E-03    |                          |                          |                           |                           |               |Jy       |2006ApJ...651...93K|no uncertainty reported|4050   A           |Broad-band measurement                                                 |043135.5 -084056 (B1950)        |Integrated from scans                                   |                                       |Averaged from previously published data                                                                                                                            
 24    |103a-O (POSS-I O)   |1.5E+01               |             |mag                 |7.40E+14 |5.77E-03    |                          |                          |                           |                           |               |Jy       |2006ApJ...651...93K|no uncertainty reported|4050   A           |Broad-band measurement                                                 |043135.5 -084056 (B1950)        |Integrated from scans                                   |                                       |Averaged from previously published data                                                                                                                            
 26    |B (OHP)             |1.6E+01               |             |mag                 |7.14E+14 |1.39E-03    |                          |                          |                           |                           |               |Jy       |1998A&AS..130..285C|no uncertainty reported|4200 A             |Broad-band measurement                                                 |04 31 35.51 -8.6783 (B1950)     |Flux integrated from map                                |Nuclear mag                            |From new raw data                                                                                                                                                  
 28    |B (B_T)             |1.4E+01               |+/-0.13      |mag                 |6.81E+14 |1.51E-02    |1.9E-03                   |1.9E-03                   |                           |                           |+/-1.91E-03    |Jy       |1991RC3.9.C...0000d|rms uncertainty        |4400       A       |Broad-band measurement                                                 |043135.5 -084042 (B1950)        |From multi-aperture data                                |                                       |Homogenized from new and previously published data; StandardJohnson UBVRI filters assumed                                                                          
 29    |B_T (VATT)          |1.4E+01               |+/-0.008     |mag                 |6.81E+14 |1.65E-02    |1.2E-04                   |1.2E-04                   |                           |                           |+/-1.22E-04    |Jy       |2005ApJ...630..784T|uncertainty            |4400   A           |Broad-band measurement                                                 |04 33 59.20 -08 35 56.3 (J2000) |Total flux                                              |                                       |From new raw data; Standard Johnson UBVRI filters assumed                                                                                                          
 30    |B (B_T^0)           |1.3E+01               |             |mag                 |6.81E+14 |2.08E-02    |                          |                          |                           |                           |               |Jy       |1991RC3.9.C...0000d|no uncertainty reported|4400       A       |Broad-band measurement                                                 |043135.5 -084042 (B1950)        |From multi-aperture data                                |                                       |Homogenized from new and previously published data;Extinction-corrected for internal and Milky Way and K-correction applied; Standard Johnson UBVRI filters assumed
 31    |g (SDSS) AB         |1.3E+01               |+/-0.05      |mag                 |6.40E+14 |2.82E-02    |1.3E-03                   |1.3E-03                   |                           |                           |+/-1.30E-03    |Jy       |2014ApJS..212...18B|uncertainty            |4681   A           |Broad-band measurement                                                 |68.50016000 -8.57923000 (J2000) |Flux in fixed aperture                                  |80"x60" aperture                       |From new raw data; Extinction-corrected for Milky Way                                                                                                              
 32    |g (SDSS) AB         |1.3E+01               |+/-0.05      |mag                 |6.40E+14 |1.70E-02    |7.8E-04                   |7.8E-04                   |                           |                           |+/-7.84E-04    |Jy       |2014ApJS..212...18B|uncertainty            |4681   A           |Broad-band measurement                                                 |68.50016000 -8.57923000 (J2000) |Flux in fixed aperture                                  |80"x60" aperture                       |From new raw data                                                                                                                                                  
 35    |V (OHP)             |1.5E+01               |             |mag                 |5.55E+14 |2.68E-03    |                          |                          |                           |                           |               |Jy       |1998A&AS..130..285C|no uncertainty reported|5400 A             |Broad-band measurement                                                 |04 31 35.51 -8.6783 (B1950)     |Flux integrated from map                                |Nuclear mag                            |From new raw data                                                                                                                                                  
 36    |V (Johnson)         |1.3E+01               |+/-0.05      |mag                 |5.42E+14 |1.62E-02    |7.6E-04                   |7.6E-04                   |                           |                           |+/-7.63E-04    |Jy       |1977ApJS...35..171H|uncertainty            |5530   A           |Broad-band measurement                                                 |                                |Flux in fixed aperture                                  |31" aperture                           |From new raw data                                                                                                                                                  
 37    |V (Johnson)         |1.4E+01               |+/-0.02      |mag                 |5.42E+14 |1.19E-02    |2.2E-04                   |2.2E-04                   |                           |                           |+/-2.22E-04    |Jy       |1979SvAL....5..305D|uncertainty            |5530   A           |Broad-band measurement                                                 |                                |Flux in fixed aperture                                  |25" aperture                           |From new raw data                                                                                                                                                  
 38    |V (Johnson)         |1.3E+01               |+/-0.05      |mag                 |5.42E+14 |1.63E-02    |7.7E-04                   |7.7E-04                   |                           |                           |+/-7.70E-04    |Jy       |1977ApJS...35..171H|uncertainty            |5530   A           |Broad-band measurement                                                 |                                |Flux in fixed aperture                                  |31" aperture                           |From new raw data                                                                                                                                                  
 39    |V (Johnson)         |1.3E+01               |+/-0.05      |mag                 |5.42E+14 |2.21E-02    |1.0E-03                   |1.0E-03                   |                           |                           |+/-1.04E-03    |Jy       |1977ApJS...35..171H|uncertainty            |5530   A           |Broad-band measurement                                                 |                                |Flux in fixed aperture                                  |43" aperture                           |From new raw data                                                                                                                                                  
 40    |V (Johnson)         |1.3E+01               |+/-0.05      |mag                 |5.42E+14 |2.17E-02    |1.0E-03                   |1.0E-03                   |                           |                           |+/-1.02E-03    |Jy       |1977ApJS...35..171H|uncertainty            |5530   A           |Broad-band measurement                                                 |                                |Flux in fixed aperture                                  |43" aperture                           |From new raw data                                                                                                                                                  
 41    |V_T (VATT)          |1.3E+01               |+/-0.013     |mag                 |5.42E+14 |2.54E-02    |3.0E-04                   |3.0E-04                   |                           |                           |+/-3.00E-04    |Jy       |2005ApJ...630..784T|uncertainty            |5530   A           |Broad-band measurement                                                 |04 33 59.20 -08 35 56.3 (J2000) |Total flux                                              |                                       |From new raw data; derived from a flux in a different bandand a color; Standard Johnson UBVRI filters assumed                                                      
 42    |V (V_T)             |1.3E+01               |+/-0.13      |mag                 |5.42E+14 |2.43E-02    |3.1E-03                   |3.1E-03                   |                           |                           |+/-3.10E-03    |Jy       |1991RC3.9.C...0000d|rms uncertainty        |5530       A       |Broad-band measurement                                                 |043135.5 -084042 (B1950)        |From multi-aperture data                                |                                       |Homogenized from new and previously published data; StandardJohnson UBVRI filters assumed                                                                          
 43    |V (V_T^0)           |1.3E+01               |             |mag                 |5.42E+14 |3.06E-02    |                          |                          |                           |                           |               |Jy       |1991RC3.9.C...0000d|no uncertainty reported|5530       A       |Broad-band measurement                                                 |043135.5 -084042 (B1950)        |From multi-aperture data                                |                                       |Homogenized from new and previously published data;Extinction-corrected for internal and Milky Way and K-correction applied; Standard Johnson UBVRI filters assumed
 44    |r (SDSS) AB         |1.2E+01               |+/-0.05      |mag                 |4.86E+14 |4.44E-02    |2.0E-03                   |2.0E-03                   |                           |                           |+/-2.04E-03    |Jy       |2014ApJS..212...18B|uncertainty            |6165   A           |Broad-band measurement                                                 |68.50016000 -8.57923000 (J2000) |Flux in fixed aperture                                  |80"x60" aperture                       |From new raw data; Extinction-corrected for Milky Way                                                                                                              
 45    |r (SDSS) AB         |1.3E+01               |+/-0.05      |mag                 |4.86E+14 |3.15E-02    |1.5E-03                   |1.5E-03                   |                           |                           |+/-1.45E-03    |Jy       |2014ApJS..212...18B|uncertainty            |6165   A           |Broad-band measurement                                                 |68.50016000 -8.57923000 (J2000) |Flux in fixed aperture                                  |80"x60" aperture                       |From new raw data                                                                                                                                                  
 54    |R (OHP)             |1.5E+01               |             |mag                 |4.41E+14 |4.44E-03    |                          |                          |                           |                           |               |Jy       |1998A&AS..130..285C|no uncertainty reported|6800 A             |Broad-band measurement                                                 |04 31 35.51 -8.6783 (B1950)     |Flux integrated from map                                |Nuclear mag                            |From new raw data                                                                                                                                                  
 55    |R_T (VATT)          |1.2E+01               |+/-0.015     |mag                 |4.33E+14 |3.76E-02    |5.2E-04                   |5.2E-04                   |                           |                           |+/-5.23E-04    |Jy       |2005ApJ...630..784T|uncertainty            |6930   A           |Broad-band measurement                                                 |04 33 59.20 -08 35 56.3 (J2000) |Total flux                                              |                                       |From new raw data; derived from a flux in a different bandand a color; Standard Johnson UBVRI filters assumed                                                      
 56    |R (Johnson)         |1.3E+01               |+/-0.02      |mag                 |4.28E+14 |2.36E-02    |4.4E-04                   |4.4E-04                   |                           |                           |+/-4.38E-04    |Jy       |1979SvAL....5..305D|uncertainty            |7000   A           |Broad-band measurement                                                 |                                |Flux in fixed aperture                                  |25" aperture                           |From new raw data; derived from a flux in a different bandand a color                                                                                              
 57    |i (SDSS) AB         |1.2E+01               |+/-0.05      |mag                 |4.01E+14 |5.48E-02    |2.5E-03                   |2.5E-03                   |                           |                           |+/-2.52E-03    |Jy       |2014ApJS..212...18B|uncertainty            |7480   A           |Broad-band measurement                                                 |68.50016000 -8.57923000 (J2000) |Flux in fixed aperture                                  |80"x60" aperture                       |From new raw data; Extinction-corrected for Milky Way                                                                                                              
 58    |i (SDSS) AB         |1.2E+01               |+/-0.05      |mag                 |4.01E+14 |4.22E-02    |1.9E-03                   |1.9E-03                   |                           |                           |+/-1.94E-03    |Jy       |2014ApJS..212...18B|uncertainty            |7480   A           |Broad-band measurement                                                 |68.50016000 -8.57923000 (J2000) |Flux in fixed aperture                                  |80"x60" aperture                       |From new raw data                                                                                                                                                  
 59    |z (SDSS) AB         |1.2E+01               |+/-0.05      |mag                 |3.36E+14 |6.73E-02    |3.1E-03                   |3.1E-03                   |                           |                           |+/-3.10E-03    |Jy       |2014ApJS..212...18B|uncertainty            |8931   A           |Broad-band measurement                                                 |68.50016000 -8.57923000 (J2000) |Flux in fixed aperture                                  |80"x60" aperture                       |From new raw data; Extinction-corrected for Milky Way                                                                                                              
 60    |z (SDSS) AB         |1.2E+01               |+/-0.05      |mag                 |3.36E+14 |5.53E-02    |2.6E-03                   |2.6E-03                   |                           |                           |+/-2.55E-03    |Jy       |2014ApJS..212...18B|uncertainty            |8931   A           |Broad-band measurement                                                 |68.50016000 -8.57923000 (J2000) |Flux in fixed aperture                                  |80"x60" aperture                       |From new raw data                                                                                                                                                  
 61    |J (UKIRT)           |3.6E+01               |+/-1.4       |milliJy             |2.50E+14 |3.58E-02    |1.4E-03                   |1.4E-03                   |                           |                           |+/-1.40E-03    |Jy       |1985ApJ...291..117L|uncertainty            |1.2 microns        |Broad-band measurement                                                 |                                |Flux in fixed aperture                                  |Aperture = 8"                          |From new raw data                                                                                                                                                  
 62    |J (KPNO)            |1.1E+01               |+/-0.05      |mag                 |2.44E+14 |4.03E-02    |1.9E-03                   |1.9E-03                   |                           |                           |+/-1.90E-03    |Jy       |1981ApJ...243..756B|uncertainty            |1.23    microns    |Broad-band measurement                                                 |                                |Flux in fixed aperture                                  |10.3" aperture                         |From new raw data                                                                                                                                                  
 63    |J (2MASS) AB        |1.2E+01               |+/-0.05      |mag                 |2.43E+14 |9.00E-02    |4.1E-03                   |4.1E-03                   |                           |                           |+/-4.14E-03    |Jy       |2014ApJS..212...18B|uncertainty            |12320   A          |Broad-band measurement                                                 |68.50016000 -8.57923000 (J2000) |Flux in fixed aperture                                  |80"x60" aperture                       |From new raw data                                                                                                                                                  
 64    |J (2MASS) AB        |1.1E+01               |+/-0.05      |mag                 |2.43E+14 |1.00E-01    |4.6E-03                   |4.6E-03                   |                           |                           |+/-4.62E-03    |Jy       |2014ApJS..212...18B|uncertainty            |12320   A          |Broad-band measurement                                                 |68.50016000 -8.57923000 (J2000) |Flux in fixed aperture                                  |80"x60" aperture                       |From new raw data; Extinction-corrected for Milky Way                                                                                                              
 65    |F_J (total)         |2.4E+00               |+/-1.85      |log milliJy         |2.41E+14 |2.75E-01    |7.1E-02                   |7.1E-02                   |                           |                           |+/-7.13E-02    |Jy       |1995ApJ...453..616S|1 sigma                |1.244      microns |Broad-band measurement                                                 |                                |Corrected to total flux from single aperture measurement|                                       |Homogenized from new and previously published data                                                                                                                 
 66    |J_14arcsec (2MASS)  |1.1E+01               |+/-0.004     |mag                 |2.40E+14 |5.02E-02    |1.9E-04                   |1.9E-04                   |                           |                           |+/-1.85E-04    |Jy       |20032MASX.C.......:|1 sigma uncert.        |1.25      microns  |Broad-band measurement                                                 |043400.03 -083444.9 (J2000)     |Flux in fixed aperture                                  |14.0 x 14.0 arcsec aperture.           |From new raw data                                                                                                                                                  
 67    |J                   |1.1E+01               |+/-0.014     |mag                 |2.40E+14 |8.95E-02    |1.2E-03                   |1.2E-03                   |                           |                           |+/-1.16E-03    |Jy       |20032MASX.C.......:|1 sigma uncert.        |1.25      microns  |Broad-band measurement                                                 |043400.03 -083444.9 (J2000)     |Flux in fixed aperture                                  |                                       |From new raw data                                                                                                                                                  
 68    |J                   |1.1E+01               |+/-0.012     |mag                 |2.40E+14 |8.02E-02    |8.9E-04                   |8.9E-04                   |                           |                           |+/-8.91E-04    |Jy       |20032MASX.C.......:|1 sigma uncert.        |1.25      microns  |Broad-band measurement                                                 |043400.03 -083444.9 (J2000)     |Flux in fixed aperture                                  |54.0 x   31.3 arcsec integration area. |From new raw data                                                                                                                                                  
 71    |F_H (total)         |2.2E+00               |+/-1.57      |log milliJy         |1.84E+14 |1.45E-01    |3.7E-02                   |3.7E-02                   |                           |                           |+/-3.74E-02    |Jy       |1995ApJ...453..616S|1 sigma                |1.634      microns |Broad-band measurement                                                 |                                |Corrected to total flux from single aperture measurement|                                       |Homogenized from new and previously published data                                                                                                                 
 73    |H_14arcsec (2MASS)  |1.0E+01               |+/-0.004     |mag                 |1.82E+14 |6.80E-02    |2.5E-04                   |2.5E-04                   |                           |                           |+/-2.51E-04    |Jy       |20032MASX.C.......:|1 sigma uncert.        |1.65      microns  |Broad-band measurement                                                 |043400.03 -083444.9 (J2000)     |Flux in fixed aperture                                  |14.0 x 14.0 arcsec aperture.           |From new raw data                                                                                                                                                  
 74    |H (UKIRT)           |5.0E+01               |+/-2.0       |milliJy             |1.82E+14 |5.00E-02    |2.0E-03                   |2.0E-03                   |                           |                           |+/-2.00E-03    |Jy       |1985ApJ...291..117L|uncertainty            |1.65 microns       |Broad-band measurement                                                 |                                |Flux in fixed aperture                                  |Aperture = 8"                          |From new raw data                                                                                                                                                  
 75    |H                   |9.9E+00               |+/-0.013     |mag                 |1.82E+14 |1.14E-01    |1.4E-03                   |1.4E-03                   |                           |                           |+/-1.37E-03    |Jy       |20032MASX.C.......:|1 sigma uncert.        |1.65      microns  |Broad-band measurement                                                 |043400.03 -083444.9 (J2000)     |Flux in fixed aperture                                  |                                       |From new raw data                                                                                                                                                  
 76    |H                   |1.0E+01               |+/-0.013     |mag                 |1.82E+14 |1.05E-01    |1.3E-03                   |1.3E-03                   |                           |                           |+/-1.26E-03    |Jy       |20032MASX.C.......:|1 sigma uncert.        |1.65      microns  |Broad-band measurement                                                 |043400.03 -083444.9 (J2000)     |Flux in fixed aperture                                  |54.0 x   31.3 arcsec integration area. |From new raw data                                                                                                                                                  
 77    |H (2MASS) AB        |1.1E+01               |+/-0.05      |mag                 |1.82E+14 |1.25E-01    |5.8E-03                   |5.8E-03                   |                           |                           |+/-5.75E-03    |Jy       |2014ApJS..212...18B|uncertainty            |16440   A          |Broad-band measurement                                                 |68.50016000 -8.57923000 (J2000) |Flux in fixed aperture                                  |80"x60" aperture                       |From new raw data; Extinction-corrected for Milky Way                                                                                                              
 78    |H (2MASS) AB        |1.1E+01               |+/-0.05      |mag                 |1.82E+14 |1.16E-01    |5.3E-03                   |5.3E-03                   |                           |                           |+/-5.34E-03    |Jy       |2014ApJS..212...18B|uncertainty            |16440   A          |Broad-band measurement                                                 |68.50016000 -8.57923000 (J2000) |Flux in fixed aperture                                  |80"x60" aperture                       |From new raw data                                                                                                                                                  
 79    |H (KPNO)            |1.1E+01               |+/-0.07      |mag                 |1.81E+14 |4.66E-02    |3.1E-03                   |3.1E-03                   |                           |                           |+/-3.10E-03    |Jy       |1981ApJ...243..756B|uncertainty            |1.66    microns    |Broad-band measurement                                                 |                                |Flux in fixed aperture                                  |10.3" aperture                         |From new raw data; derived from a flux in a different bandand a color                                                                                              
 84    |Ks (2MASS) AB       |1.1E+01               |+/-0.05      |mag                 |1.39E+14 |1.17E-01    |5.4E-03                   |5.4E-03                   |                           |                           |+/-5.40E-03    |Jy       |2014ApJS..212...18B|uncertainty            |21590   A          |Broad-band measurement                                                 |68.50016000 -8.57923000 (J2000) |Flux in fixed aperture                                  |80"x60" aperture                       |From new raw data; Extinction-corrected for Milky Way                                                                                                              
 85    |Ks (2MASS) AB       |1.1E+01               |+/-0.05      |mag                 |1.39E+14 |1.12E-01    |5.1E-03                   |5.1E-03                   |                           |                           |+/-5.14E-03    |Jy       |2014ApJS..212...18B|uncertainty            |21590   A          |Broad-band measurement                                                 |68.50016000 -8.57923000 (J2000) |Flux in fixed aperture                                  |80"x60" aperture                       |From new raw data                                                                                                                                                  
 86    |K_s                 |9.5E+00               |+/-0.020     |mag                 |1.38E+14 |1.09E-01    |2.0E-03                   |2.0E-03                   |                           |                           |+/-2.02E-03    |Jy       |20032MASX.C.......:|1 sigma uncert.        |2.17      microns  |Broad-band measurement                                                 |043400.03 -083444.9 (J2000)     |Flux in fixed aperture                                  |                                       |From new raw data                                                                                                                                                  
 87    |K_s_14arcsec (2MASS)|9.9E+00               |+/-0.005     |mag                 |1.38E+14 |7.05E-02    |3.3E-04                   |3.3E-04                   |                           |                           |+/-3.26E-04    |Jy       |20032MASX.C.......:|1 sigma uncert.        |2.17      microns  |Broad-band measurement                                                 |043400.03 -083444.9 (J2000)     |Flux in fixed aperture                                  |14.0 x 14.0 arcsec aperture.           |From new raw data                                                                                                                                                  
 88    |K_s                 |9.5E+00               |+/-0.020     |mag                 |1.38E+14 |1.01E-01    |1.9E-03                   |1.9E-03                   |                           |                           |+/-1.89E-03    |Jy       |20032MASX.C.......:|1 sigma uncert.        |2.17      microns  |Broad-band measurement                                                 |043400.03 -083444.9 (J2000)     |Flux in fixed aperture                                  |54.0 x   31.3 arcsec integration area. |From new raw data                                                                                                                                                  
 90    |F_K (total)         |2.1E+00               |+/-1.46      |log milliJy         |1.37E+14 |1.12E-01    |2.9E-02                   |2.9E-02                   |                           |                           |+/-2.91E-02    |Jy       |1995ApJ...453..616S|1 sigma                |2.194      microns |Broad-band measurement                                                 |                                |Corrected to total flux from single aperture measurement|                                       |Homogenized from new and previously published data                                                                                                                 
 91    |K (UKIRT)           |5.1E+01               |+/-2.0       |milliJy             |1.36E+14 |5.11E-02    |2.0E-03                   |2.0E-03                   |                           |                           |+/-2.00E-03    |Jy       |1985ApJ...291..117L|uncertainty            |2.2 microns        |Broad-band measurement                                                 |                                |Flux in fixed aperture                                  |Aperture = 8"                          |From new raw data                                                                                                                                                  
 92    |K (KPNO)            |1.0E+01               |+/-0.10      |mag                 |1.35E+14 |5.32E-02    |5.1E-03                   |5.1E-03                   |                           |                           |+/-5.13E-03    |Jy       |1981ApJ...243..756B|uncertainty            |2.22    microns    |Broad-band measurement                                                 |                                |Flux in fixed aperture                                  |10.3" aperture                         |From new raw data; derived from a flux in a different bandand a color                                                                                              
 97    |3.4 microns WISE AB |1.2E+01               |+/-0.10      |mag                 |8.93E+13 |8.80E-02    |8.1E-03                   |8.1E-03                   |                           |                           |+/-8.11E-03    |Jy       |2014ApJS..212...18B|uncertainty            |33570   A          |Broad-band measurement                                                 |68.50016000 -8.57923000 (J2000) |Flux in fixed aperture                                  |80"x60" aperture                       |From new raw data; Extinction-corrected for Milky Way                                                                                                              
 98    |3.4 microns WISE AB |1.2E+01               |+/-0.10      |mag                 |8.93E+13 |8.56E-02    |7.9E-03                   |7.9E-03                   |                           |                           |+/-7.88E-03    |Jy       |2014ApJS..212...18B|uncertainty            |33570   A          |Broad-band measurement                                                 |68.50016000 -8.57923000 (J2000) |Flux in fixed aperture                                  |80"x60" aperture                       |From new raw data                                                                                                                                                  
 99    |L (UKIRT)           |6.5E+01               |+/-2.6       |milliJy             |8.57E+13 |6.53E-02    |2.6E-03                   |2.6E-03                   |                           |                           |+/-2.60E-03    |Jy       |1985ApJ...291..117L|uncertainty            |3.5 microns        |Broad-band measurement                                                 |                                |Flux in fixed aperture                                  |Aperture = 8"                          |From new raw data                                                                                                                                                  
 100   |L (UKIRT)           |5.8E+01               |+/-3.1       |milliJy             |8.57E+13 |5.80E-02    |3.1E-03                   |3.1E-03                   |                           |                           |+/-3.10E-03    |Jy       |1985ApJ...291..117L|uncertainty            |3.5 microns        |Broad-band measurement                                                 |                                |Flux in fixed aperture                                  |Aperture = 5"                          |From new raw data                                                                                                                                                  
 101   |3.6 microns IRAC AB |1.1E+01               |+/-0.10      |mag                 |8.46E+13 |9.43E-02    |8.7E-03                   |8.7E-03                   |                           |                           |+/-8.69E-03    |Jy       |2014ApJS..212...18B|uncertainty            |35440   A          |Broad-band measurement                                                 |68.50016000 -8.57923000 (J2000) |Flux in fixed aperture                                  |80"x60" aperture                       |From new raw data                                                                                                                                                  
 102   |3.6 microns IRAC AB |1.1E+01               |+/-0.10      |mag                 |8.46E+13 |9.68E-02    |8.9E-03                   |8.9E-03                   |                           |                           |+/-8.92E-03    |Jy       |2014ApJS..212...18B|uncertainty            |35440   A          |Broad-band measurement                                                 |68.50016000 -8.57923000 (J2000) |Flux in fixed aperture                                  |80"x60" aperture                       |From new raw data; Extinction-corrected for Milky Way                                                                                                              
 103   |3.6 microns (IRAC)  |1.0E-01               |+/-3.09E-3   |Jy                  |8.44E+13 |1.03E-01    |3.1E-03                   |3.1E-03                   |                           |                           |+/-3.09E-03    |Jy       |2008ApJ...678..804E|rms uncertainty        |3.550 microns      |Broad-band measurement                                                 |04 34 00.1 -08 34 44.9 (J2000)  |Corrected to total flux from single aperture measurement|Color-corrected                        |From new raw data                                                                                                                                                  
 105   |4.5 microns IRAC AB |1.2E+01               |+/-0.10      |mag                 |6.68E+13 |7.91E-02    |7.3E-03                   |7.3E-03                   |                           |                           |+/-7.28E-03    |Jy       |2014ApJS..212...18B|uncertainty            |44870   A          |Broad-band measurement                                                 |68.50016000 -8.57923000 (J2000) |Flux in fixed aperture                                  |80"x60" aperture                       |From new raw data; Extinction-corrected for Milky Way                                                                                                              
 106   |4.5 microns IRAC AB |1.2E+01               |+/-0.10      |mag                 |6.68E+13 |7.74E-02    |7.1E-03                   |7.1E-03                   |                           |                           |+/-7.13E-03    |Jy       |2014ApJS..212...18B|uncertainty            |44870   A          |Broad-band measurement                                                 |68.50016000 -8.57923000 (J2000) |Flux in fixed aperture                                  |80"x60" aperture                       |From new raw data                                                                                                                                                  
 107   |4.5 microns (IRAC)  |7.6E-02               |+/-2.27E-3   |Jy                  |6.67E+13 |7.56E-02    |2.3E-03                   |2.3E-03                   |                           |                           |+/-2.27E-03    |Jy       |2008ApJ...678..804E|rms uncertainty        |4.493 microns      |Broad-band measurement                                                 |04 34 00.1 -08 34 44.9 (J2000)  |Corrected to total flux from single aperture measurement|Color-corrected                        |From new raw data                                                                                                                                                  
 108   |4.6 microns WISE AB |1.2E+01               |+/-0.10      |mag                 |6.51E+13 |7.40E-02    |6.8E-03                   |6.8E-03                   |                           |                           |+/-6.81E-03    |Jy       |2014ApJS..212...18B|uncertainty            |46060   A          |Broad-band measurement                                                 |68.50016000 -8.57923000 (J2000) |Flux in fixed aperture                                  |80"x60" aperture                       |From new raw data; Extinction-corrected for Milky Way                                                                                                              
 109   |4.6 microns WISE AB |1.2E+01               |+/-0.10      |mag                 |6.51E+13 |7.25E-02    |6.7E-03                   |6.7E-03                   |                           |                           |+/-6.68E-03    |Jy       |2014ApJS..212...18B|uncertainty            |46060   A          |Broad-band measurement                                                 |68.50016000 -8.57923000 (J2000) |Flux in fixed aperture                                  |80"x60" aperture                       |From new raw data                                                                                                                                                  
 110   |M (UKIRT)           |4.8E+01               |+/-10.1      |milliJy             |6.25E+13 |4.75E-02    |1.0E-02                   |1.0E-02                   |                           |                           |+/-1.01E-02    |Jy       |1985ApJ...291..117L|uncertainty            |4.8 microns        |Broad-band measurement                                                 |                                |Flux in fixed aperture                                  |Aperture = 5"                          |From new raw data                                                                                                                                                  
 111   |5.0 microns         |9.2E-01               |+/-0.05      |Jy                  |6.00E+13 |9.20E-01    |5.0E-02                   |5.0E-02                   |                           |                           |+/-5.00E-02    |Jy       |1972ApJ...176L..95R|1 sigma                |5.0 microns        |Broad-band measurement                                                 |                                |Flux in fixed aperture                                  |6" aperture                            |From new raw data                                                                                                                                                  
 112   |5.0 microns         |1.0E+00               |+/-0.11      |Jy                  |6.00E+13 |2.70E-01    |1.1E-01                   |1.1E-01                   |                           |                           |+/-1.10E-01    |Jy       |1972ApJ...176L..95R|1 sigma                |5.0 microns        |Broad-band measurement                                                 |                                |Flux in fixed aperture                                  |6" aperture                            |From new raw data                                                                                                                                                  
 114   |5.8 microns IRAC AB |1.0E+01               |+/-0.10      |mag                 |5.25E+13 |2.89E-01    |2.7E-02                   |2.7E-02                   |                           |                           |+/-2.66E-02    |Jy       |2014ApJS..212...18B|uncertainty            |57100   A          |Broad-band measurement                                                 |68.50016000 -8.57923000 (J2000) |Flux in fixed aperture                                  |80"x60" aperture                       |From new raw data                                                                                                                                                  
 115   |5.8 microns IRAC AB |1.0E+01               |+/-0.10      |mag                 |5.25E+13 |2.93E-01    |2.7E-02                   |2.7E-02                   |                           |                           |+/-2.70E-02    |Jy       |2014ApJS..212...18B|uncertainty            |57100   A          |Broad-band measurement                                                 |68.50016000 -8.57923000 (J2000) |Flux in fixed aperture                                  |80"x60" aperture                       |From new raw data; Extinction-corrected for Milky Way                                                                                                              
 116   |5.8 microns (IRAC)  |2.9E-01               |+/-8.81E-3   |Jy                  |5.23E+13 |2.93E-01    |8.8E-03                   |8.8E-03                   |                           |                           |+/-8.81E-03    |Jy       |2008ApJ...678..804E|rms uncertainty        |5.731 microns      |Broad-band measurement                                                 |04 34 00.1 -08 34 44.9 (J2000)  |Corrected to total flux from single aperture measurement|Color-corrected                        |From new raw data                                                                                                                                                  
 117   |6 microns (IRS)     |1.4E-01               |             |Jy                  |5.00E+13 |1.40E-01    |                          |                          |                           |                           |               |Jy       |2006ApJ...653.1129B|no uncertainty reported|6   microns        |Broad-band measurement                                                 |04 33 59.85 -08 34 44.0 (J2000) |Flux integrated from map                                |                                       |From new raw data                                                                                                                                                  
 122   |8.0 microns (IRAC)  |8.9E-01               |+/-2.66E-2   |Jy                  |3.81E+13 |8.87E-01    |2.7E-02                   |2.7E-02                   |                           |                           |+/-2.66E-02    |Jy       |2008ApJ...678..804E|rms uncertainty        |7.872 microns      |Broad-band measurement                                                 |04 34 00.1 -08 34 44.9 (J2000)  |Corrected to total flux from single aperture measurement|Color-corrected                        |From new raw data                                                                                                                                                  
 125   |Si2 (GeminiS)       |                      |<420.3       |milliJy             |3.43E+13 |            |                          |                          |4.2E-01                    |                           |<4.20E-01      |Jy       |2014MNRAS.439.1648A|3 sigma                |8.74   microns     |Broad-band measurement                                                 |068.499583 -08.578889 (J2000)   |Flux in fixed aperture                                  |Nuclear flux                           |From reprocessed raw data                                                                                                                                          
 126   |Si2 (GeminiS)       |                      |<397.7       |milliJy             |3.43E+13 |            |                          |                          |4.0E-01                    |                           |<3.98E-01      |Jy       |2014MNRAS.439.1648A|3 sigma                |8.74   microns     |Broad-band measurement                                                 |068.499583 -08.578889 (J2000)   |Flux in fixed aperture                                  |Nuclear flux                           |From reprocessed raw data                                                                                                                                          
 127   |10.5 microns        |1.0E+00               |+/-0.03      |Jy                  |2.86E+13 |1.02E+00    |3.0E-02                   |3.0E-02                   |                           |                           |+/-3.00E-02    |Jy       |1972ApJ...176L..95R|1 sigma                |10.5 microns       |Broad-band measurement                                                 |                                |Flux in fixed aperture                                  |6" aperture                            |From new raw data                                                                                                                                                  
 128   |10.6 microns        |6.3E-01               |             |Jy                  |2.83E+13 |6.30E-01    |                          |                          |                           |                           |               |Jy       |1979ApJ...229..111L|no uncertainty reported|10.6     microns   |Broad-band measurement                                                 |                                |Flux in fixed aperture                                  |8.5" aperture                          |From new raw data                                                                                                                                                  
 129   |PAH2 11.25 (VLT)    |7.2E+02               |             |milliJy             |2.66E+13 |7.20E-01    |                          |                          |                           |                           |               |Jy       |2008A&A...488...83S|no uncertainty reported|11.25 microns      |Broad-band measurement                                                 |                                |Flux integrated from map                                |                                       |From new raw data                                                                                                                                                  
 130   |PAH2 (VLT)          |                      |<731.4       |milliJy             |2.66E+13 |            |                          |                          |7.3E-01                    |                           |<7.31E-01      |Jy       |2014MNRAS.439.1648A|3 sigma                |11.25   microns    |Broad-band measurement                                                 |068.499583 -08.578889 (J2000)   |Flux in fixed aperture                                  |Nuclear flux                           |From reprocessed raw data                                                                                                                                          
 133   |11.7 microns        |1.0E+03               |+/-103       |milliJy             |2.56E+13 |1.03E+00    |1.0E-01                   |1.0E-01                   |                           |                           |+/-1.03E-01    |Jy       |2001AJ....122.1213S|estimated error        |11.7       microns |Broad-band measurement                                                 |                                |Flux in fixed aperture                                  |4" aperture                            |From new raw data                                                                                                                                                  
 134   |12 microns WISE AB  |8.7E+00               |+/-0.10      |mag                 |2.54E+13 |1.21E+00    |1.1E-01                   |1.1E-01                   |                           |                           |+/-1.11E-01    |Jy       |2014ApJS..212...18B|uncertainty            |118100   A         |Broad-band measurement                                                 |68.50016000 -8.57923000 (J2000) |Flux in fixed aperture                                  |80"x60" aperture                       |From new raw data                                                                                                                                                  
 135   |12 microns WISE AB  |8.7E+00               |+/-0.10      |mag                 |2.54E+13 |1.22E+00    |1.1E-01                   |1.1E-01                   |                           |                           |+/-1.12E-01    |Jy       |2014ApJS..212...18B|uncertainty            |118100   A         |Broad-band measurement                                                 |68.50016000 -8.57923000 (J2000) |Flux in fixed aperture                                  |80"x60" aperture                       |From new raw data; Extinction-corrected for Milky Way                                                                                                              
 136   |12 microns (IRAS)   |1.4E+00               |+/-0.023     |Jy                  |2.50E+13 |1.38E+00    |2.3E-02                   |2.3E-02                   |                           |                           |+/-2.30E-02    |Jy       |2003AJ....126.1607S|1 sigma                |12   microns       |Broad-band measurement                                                 |04 34 00.1 -08 34 46 (J2000)    |Total flux                                              |Size, Method, Flag codes: UT;see paper |From reprocessed raw data                                                                                                                                          
 137   |12 microns (IRAS)   |1.4E+00               |+/-0.033     |Jy                  |2.50E+13 |1.44E+00    |3.3E-02                   |3.3E-02                   |                           |                           |+/-3.30E-02    |Jy       |1989AJ.....98..766S|rms noise              |12         microns |Broad-band measurement                                                 |043135.8 -084055 (B1950)        |Integrated from scans                                   |Unresolved with 0.77' beam             |From reprocessed raw data                                                                                                                                          
 138   |12 microns (IRAS)   |1.4E+00               |+/-5   %     |Jy                  |2.50E+13 |1.44E+00    |7.2E-02                   |7.2E-02                   |                           |                           |+/-7.21E-02    |Jy       |1990IRASF.C...0000M|uncertainty            |12        microns  |Broad-band measurement                                                 |043135.8 -084058 (B1950)        |Flux in fixed aperture                                  |IRAS quality flag = 3                  |From new raw data                                                                                                                                                  
 139   |12.5 microns        |1.2E+03               |+/-122       |milliJy             |2.40E+13 |1.22E+00    |1.2E-01                   |1.2E-01                   |                           |                           |+/-1.22E-01    |Jy       |2001AJ....122.1213S|estimated error        |12.5       microns |Broad-band measurement                                                 |                                |Flux in fixed aperture                                  |4" aperture                            |From new raw data                                                                                                                                                  
 144   |15 microns (IRS)    |1.1E+00               |             |Jy                  |2.00E+13 |1.10E+00    |                          |                          |                           |                           |               |Jy       |2006ApJ...653.1129B|no uncertainty reported|15   microns       |Broad-band measurement                                                 |04 33 59.85 -08 34 44.0 (J2000) |Flux integrated from map                                |                                       |From new raw data                                                                                                                                                  
 148   |17.7 microns Subaru |3.0E+03               |             |milliJy             |1.69E+13 |2.97E+00    |                          |                          |                           |                           |               |Jy       |2011AJ....141..156I|no uncertainty reported|17.7 microns       |Broad-band measurement                                                 |                                |Flux in fixed aperture                                  |                                       |From new raw data                                                                                                                                                  
 149   |Q17.7 (Subaru)      |                      |<2572.9      |milliJy             |1.69E+13 |            |                          |                          |2.6E+00                    |                           |<2.57E+00      |Jy       |2014MNRAS.439.1648A|3 sigma                |17.69   microns    |Broad-band measurement                                                 |068.499583 -08.578889 (J2000)   |Flux in fixed aperture                                  |Nuclear flux                           |From reprocessed raw data                                                                                                                                          
 152   |Q2 (VLT)            |                      |<2666.3      |milliJy             |1.60E+13 |            |                          |                          |2.7E+00                    |                           |<2.67E+00      |Jy       |2014MNRAS.439.1648A|3 sigma                |18.72   microns    |Broad-band measurement                                                 |068.499583 -08.578889 (J2000)   |Flux in fixed aperture                                  |Nuclear flux                           |From reprocessed raw data                                                                                                                                          
 153   |21 microns          |1.0E+00               |+/-0.3       |Jy                  |1.43E+13 |4.00E+00    |3.0E-01                   |3.0E-01                   |                           |                           |+/-3.00E-01    |Jy       |1972ApJ...176L..95R|1 sigma                |21 microns         |Broad-band measurement                                                 |                                |Flux in fixed aperture                                  |6" aperture                            |From new raw data                                                                                                                                                  
 154   |21 microns          |3.1E+00               |+/-0.3       |Jy                  |1.43E+13 |3.10E+00    |3.0E-01                   |3.0E-01                   |                           |                           |+/-3.00E-01    |Jy       |1979ApJ...229..111L|uncertainty            |21       microns   |Broad-band measurement                                                 |                                |Flux in fixed aperture                                  |8.5" aperture                          |Recalibrated data                                                                                                                                                  
 155   |22 microns WISE AB  |7.1E+00               |+/-0.10      |mag                 |1.35E+13 |5.49E+00    |5.1E-01                   |5.1E-01                   |                           |                           |+/-5.05E-01    |Jy       |2014ApJS..212...18B|uncertainty            |221400   A         |Broad-band measurement                                                 |68.50016000 -8.57923000 (J2000) |Flux in fixed aperture                                  |80"x60" aper; Filter curve corr        |From new raw data; Extinction-corrected for Milky Way                                                                                                              
 156   |22 microns WISE AB  |7.1E+00               |+/-0.10      |mag                 |1.35E+13 |5.46E+00    |5.0E-01                   |5.0E-01                   |                           |                           |+/-5.03E-01    |Jy       |2014ApJS..212...18B|uncertainty            |221400   A         |Broad-band measurement                                                 |68.50016000 -8.57923000 (J2000) |Flux in fixed aperture                                  |80"x60" aper; Filter curve corr        |From new raw data                                                                                                                                                  
 157   |22 microns WISE AB  |6.9E+00               |+/-0.10      |mag                 |1.35E+13 |6.31E+00    |5.8E-01                   |5.8E-01                   |                           |                           |+/-5.81E-01    |Jy       |2014ApJS..212...18B|uncertainty            |221400   A         |Broad-band measurement                                                 |68.50016000 -8.57923000 (J2000) |Flux in fixed aperture                                  |80"x60" aperture                       |From new raw data                                                                                                                                                  
 158   |22 microns WISE AB  |6.9E+00               |+/-0.10      |mag                 |1.35E+13 |6.34E+00    |5.8E-01                   |5.8E-01                   |                           |                           |+/-5.84E-01    |Jy       |2014ApJS..212...18B|uncertainty            |221400   A         |Broad-band measurement                                                 |68.50016000 -8.57923000 (J2000) |Flux in fixed aperture                                  |80"x60" aperture                       |From new raw data; Extinction-corrected for Milky Way                                                                                                              
 159   |24 microns MIPS AB  |7.0E+00               |+/-0.10      |mag                 |1.28E+13 |5.88E+00    |5.4E-01                   |5.4E-01                   |                           |                           |+/-5.41E-01    |Jy       |2014ApJS..212...18B|uncertainty            |235100   A         |Broad-band measurement                                                 |68.50016000 -8.57923000 (J2000) |Flux in fixed aperture                                  |80"x60" aperture                       |From new raw data; Extinction-corrected for Milky Way                                                                                                              
 160   |24 microns MIPS AB  |7.0E+00               |+/-0.10      |mag                 |1.28E+13 |5.85E+00    |5.4E-01                   |5.4E-01                   |                           |                           |+/-5.39E-01    |Jy       |2014ApJS..212...18B|uncertainty            |235100   A         |Broad-band measurement                                                 |68.50016000 -8.57923000 (J2000) |Flux in fixed aperture                                  |80"x60" aperture                       |From new raw data                                                                                                                                                  
 161   |24 microns (MIPS)   |5.9E+00               |+/-1.18E-1   |Jy                  |1.27E+13 |5.89E+00    |1.2E-01                   |1.2E-01                   |                           |                           |+/-1.18E-01    |Jy       |2008ApJ...678..804E|rms uncertainty        |23.68 microns      |Broad-band measurement                                                 |04 34 00.1 -08 34 44.9 (J2000)  |Corrected to total flux from single aperture measurement|Color-corrected                        |From new raw data                                                                                                                                                  
 163   |24.5 microns        |7.0E+00               |+/-0.7       |Jy                  |1.22E+13 |7.00E+00    |7.0E-01                   |7.0E-01                   |                           |                           |+/-7.00E-01    |Jy       |2001AJ....122.1213S|estimated error        |24.5       microns |Broad-band measurement                                                 |                                |Flux in fixed aperture                                  |4" aperture                            |From new raw data                                                                                                                                                  
 164   |25 microns (IRAS)   |7.5E+00               |+/-0.025     |Jy                  |1.20E+13 |7.50E+00    |2.5E-02                   |2.5E-02                   |                           |                           |+/-2.50E-02    |Jy       |2003AJ....126.1607S|1 sigma                |25   microns       |Broad-band measurement                                                 |04 34 00.1 -08 34 46 (J2000)    |Total flux                                              |Size, Method, Flag codes: UT;see paper |From reprocessed raw data                                                                                                                                          
 165   |25 microns (IRAS)   |7.3E+00               |+/-5   %     |Jy                  |1.20E+13 |7.29E+00    |7.2E-02                   |7.2E-02                   |                           |                           |+/-7.21E-02    |Jy       |1990IRASF.C...0000M|uncertainty            |25        microns  |Broad-band measurement                                                 |043135.8 -084058 (B1950)        |Flux in fixed aperture                                  |IRAS quality flag = 3                  |From new raw data                                                                                                                                                  
 166   |25 microns (IRAS)   |7.8E+00               |+/-0.028     |Jy                  |1.20E+13 |7.82E+00    |2.8E-02                   |2.8E-02                   |                           |                           |+/-2.80E-02    |Jy       |1989AJ.....98..766S|rms noise              |25         microns |Broad-band measurement                                                 |043135.8 -084055 (B1950)        |Integrated from scans                                   |Unresolved with 0.78' beam             |From reprocessed raw data                                                                                                                                          
 169   |30 microns (IRS)    |5.8E+00               |             |Jy                  |9.99E+12 |5.80E+00    |                          |                          |                           |                           |               |Jy       |2006ApJ...653.1129B|no uncertainty reported|30   microns       |Broad-band measurement                                                 |04 33 59.85 -08 34 44.0 (J2000) |Flux integrated from map                                |                                       |From new raw data                                                                                                                                                  
 174   |52 microns (ISO)    |2.6E+01               |+/-2.6       |Jy                  |5.77E+12 |2.56E+01    |2.6E+00                   |2.6E+00                   |                           |                           |+/-2.60E+00    |Jy       |2008ApJS..178..280B|uncertainty            |52 microns         |Broad-band measurement                                                 |04 34 00.03 -08 34 43.7 (J2000) |Flux integrated from map                                |                                       |From new raw data                                                                                                                                                  
 175   |57 microns (ISO)    |3.1E+01               |+/-3.0       |Jy                  |5.26E+12 |3.07E+01    |3.0E+00                   |3.0E+00                   |                           |                           |+/-3.00E+00    |Jy       |2008ApJS..178..280B|uncertainty            |57 microns         |Broad-band measurement                                                 |04 34 00.03 -08 34 43.7 (J2000) |Flux integrated from map                                |                                       |From new raw data                                                                                                                                                  
 176   |60 microns (IRAS)   |3.2E+01               |+/-0.083     |Jy                  |5.00E+12 |3.21E+01    |8.3E-02                   |8.3E-02                   |                           |                           |+/-8.30E-02    |Jy       |2003AJ....126.1607S|1 sigma                |60   microns       |Broad-band measurement                                                 |04 34 00.1 -08 34 46 (J2000)    |Total flux                                              |Size, Method, Flag codes: UT;see paper |From reprocessed raw data                                                                                                                                          
 177   |60 microns (IRAS)   |3.3E+01               |+/-0.093     |Jy                  |5.00E+12 |3.31E+01    |9.3E-02                   |9.3E-02                   |                           |                           |+/-9.30E-02    |Jy       |1989AJ.....98..766S|rms noise              |60         microns |Broad-band measurement                                                 |043135.8 -084055 (B1950)        |Integrated from scans                                   |Unresolved with 1.44' beam             |From reprocessed raw data                                                                                                                                          
 178   |60 microns (IRAS)   |3.2E+01               |+/-4   %     |Jy                  |5.00E+12 |3.23E+01    |1.3E+00                   |1.3E+00                   |                           |                           |+/-1.29E+00    |Jy       |1990IRASF.C...0000M|uncertainty            |60        microns  |Broad-band measurement                                                 |043135.8 -084058 (B1950)        |Flux in fixed aperture                                  |IRAS quality flag = 2                  |From new raw data                                                                                                                                                  
 179   |63 microns (ISO)    |4.3E+01               |+/-4.4       |Jy                  |4.76E+12 |4.31E+01    |4.4E+00                   |4.4E+00                   |                           |                           |+/-4.40E+00    |Jy       |2008ApJS..178..280B|uncertainty            |63 microns         |Broad-band measurement                                                 |04 34 00.03 -08 34 43.7 (J2000) |Flux integrated from map                                |                                       |From new raw data                                                                                                                                                  
 181   |70 microns (MIPS)   |2.5E+01               |+/-1.24E+0   |Jy                  |4.20E+12 |2.48E+01    |1.2E+00                   |1.2E+00                   |                           |                           |+/-1.24E+00    |Jy       |2008ApJ...678..804E|rms uncertainty        |71.42 microns      |Broad-band measurement                                                 |04 34 00.1 -08 34 44.9 (J2000)  |Corrected to total flux from single aperture measurement|Color-corrected                        |From new raw data                                                                                                                                                  
 182   |88 microns (ISO)    |4.9E+01               |+/-4.9       |Jy                  |3.41E+12 |4.92E+01    |4.9E+00                   |4.9E+00                   |                           |                           |+/-4.90E+00    |Jy       |2008ApJS..178..280B|uncertainty            |88 microns         |Broad-band measurement                                                 |04 34 00.03 -08 34 43.7 (J2000) |Flux integrated from map                                |                                       |From new raw data                                                                                                                                                  
 183   |100 microns (IRAS)  |3.4E+01               |+/-0.43      |Jy                  |3.00E+12 |3.43E+01    |4.3E-01                   |4.3E-01                   |                           |                           |+/-4.30E-01    |Jy       |2003AJ....126.1607S|1 sigma                |100   microns      |Broad-band measurement                                                 |04 34 00.1 -08 34 46 (J2000)    |Total flux                                              |Size, Method, Flag codes: UT;see paper |From reprocessed raw data                                                                                                                                          
 184   |100 microns (IRAS)  |3.6E+01               |+/-0.48      |Jy                  |3.00E+12 |3.62E+01    |4.8E-01                   |4.8E-01                   |                           |                           |+/-4.80E-01    |Jy       |1989AJ.....98..766S|rms noise              |100        microns |Broad-band measurement                                                 |043135.8 -084055 (B1950)        |Integrated from scans                                   |Unresolved with 2.94' beam             |From reprocessed raw data                                                                                                                                          
 185   |100 microns (IRAS)  |3.3E+01               |+/-4   %     |Jy                  |3.00E+12 |3.27E+01    |1.3E+00                   |1.3E+00                   |                           |                           |+/-1.31E+00    |Jy       |1990IRASF.C...0000M|uncertainty            |100       microns  |Broad-band measurement                                                 |043135.8 -084058 (B1950)        |Flux in fixed aperture                                  |IRAS quality flag = 2                  |From new raw data                                                                                                                                                  
 186   |122 microns (ISO)   |2.5E+01               |+/-2.1       |Jy                  |2.46E+12 |2.50E+01    |2.1E+00                   |2.1E+00                   |                           |                           |+/-2.10E+00    |Jy       |2008ApJS..178..280B|uncertainty            |122 microns        |Broad-band measurement                                                 |04 34 00.03 -08 34 43.7 (J2000) |Flux integrated from map                                |                                       |From new raw data                                                                                                                                                  
 188   |145 microns (ISO)   |2.0E+01               |+/-1.9       |Jy                  |2.07E+12 |2.03E+01    |1.9E+00                   |1.9E+00                   |                           |                           |+/-1.90E+00    |Jy       |2008ApJS..178..280B|uncertainty            |145 microns        |Broad-band measurement                                                 |04 34 00.03 -08 34 43.7 (J2000) |Flux integrated from map                                |                                       |From new raw data                                                                                                                                                  
 189   |160 microns (MIPS)  |1.7E+01               |+/-2.05E+0   |Jy                  |1.92E+12 |1.71E+01    |2.1E+00                   |2.1E+00                   |                           |                           |+/-2.05E+00    |Jy       |2008ApJ...678..804E|rms uncertainty        |155.90 microns     |Broad-band measurement                                                 |04 34 00.1 -08 34 44.9 (J2000)  |Corrected to total flux from single aperture measurement|Color-corrected                        |From new raw data                                                                                                                                                  
 190   |158 microns (ISO)   |1.6E+01               |+/-2.2       |Jy                  |1.90E+12 |1.63E+01    |2.2E+00                   |2.2E+00                   |                           |                           |+/-2.20E+00    |Jy       |2008ApJS..178..280B|uncertainty            |158 microns        |Broad-band measurement                                                 |04 34 00.03 -08 34 43.7 (J2000) |Flux integrated from map                                |                                       |From new raw data                                                                                                                                                  
 192   |170 microns (ISO)   |1.3E+01               |+/-1.2       |Jy                  |1.76E+12 |1.25E+01    |1.2E+00                   |1.2E+00                   |                           |                           |+/-1.20E+00    |Jy       |2008ApJS..178..280B|uncertainty            |170 microns        |Broad-band measurement                                                 |04 34 00.03 -08 34 43.7 (J2000) |Flux integrated from map                                |                                       |From new raw data                                                                                                                                                  
 193   |170 microns (ISO)   |1.6E+01               |+/-15  %     |Jy                  |1.76E+12 |1.63E+01    |2.4E+00                   |2.4E+00                   |                           |                           |+/-2.44E+00    |Jy       |2004A&A...422...39S|uncertainty            |170      microns   |Broad-band measurement                                                 |04 34 00.14 -08 34 57.1 (J2000) |Integrated from scans                                   |                                       |Averaged from previously published data                                                                                                                            
 194   |350 microns (CSO)   |1.2E+00               |+/-0.05      |Jy                  |8.57E+11 |1.18E+00    |5.0E-02                   |5.0E-02                   |                           |                           |+/-5.00E-02    |Jy       |2007ApJ...662..284Y|uncertainty            |350   microns      |Broad-band measurement                                                 |04 33 59.8 -08 34 44 (J2000)    |Flux integrated from map                                |                                       |From new raw data                                                                                                                                                  
 195   |350 microns         |                      |<3.2         |Jy                  |8.57E+11 |            |                          |                          |3.2E+00                    |                           |<3.20E+00      |Jy       |1989ApJ...339..859E|3 sigma                |350   microns      |Broad-band measurement                                                 |                                |Flux in fixed aperture                                  |104" aperture                          |From new raw data                                                                                                                                                  
 196   |350 microns         |1.9E+00               |+/-0.43      |Jy                  |8.57E+11 |1.87E+00    |4.3E-01                   |4.3E-01                   |                           |                           |+/-4.30E-01    |Jy       |1999CIT...T00R....B|1 sigma                |350        microns |Broad-band measurement                                                 |                                |Flux integrated from map                                |                                       |From new raw data                                                                                                                                                  
 197   |450 microns (SCUBA) |9.8E+02               |+/-167       |milliJy             |6.66E+11 |9.81E-01    |1.7E-01                   |1.7E-01                   |                           |                           |+/-1.67E-01    |Jy       |2001MNRAS.327..697D|uncertainty            |450   microns      |Broad-band measurement                                                 |04 34 00.0 -08 34 45 (J2000)    |Modelled datum; Beam filling or dilution corrected      |                                       |Averaged new and previously published data                                                                                                                         
 201   |850 microns (SCUBA) |2.2E+02               |+/-32        |milliJy             |3.53E+11 |2.19E-01    |3.2E-02                   |3.2E-02                   |                           |                           |+/-3.20E-02    |Jy       |2000MNRAS.315..115D|uncertainty            |850       microns  |Broad-band measurement                                                 |043400.0 -083445 (J2000)        |Flux integrated from map                                |                                       |From new raw data; Corrected for contaminating sources                                                                                                             
 202   |880 microns (SMA)   |2.7E+01               |+/-7         |milliJy             |3.41E+11 |2.70E-02    |7.0E-03                   |7.0E-03                   |                           |                           |+/-7.00E-03    |Jy       |2008ApJS..178..189W|uncertainty            |880 microns        |Broad-band measurement                                                 |                                |Flux integrated from map                                |                                       |From new raw data                                                                                                                                                  
 203   |1.3 mm (SMA)        |2.1E+01               |+/-3         |milliJy             |2.31E+11 |2.10E-02    |3.0E-03                   |3.0E-03                   |                           |                           |+/-3.00E-03    |Jy       |2008ApJS..178..189W|uncertainty            |1.3 mm             |Broad-band measurement                                                 |                                |Flux integrated from map                                |                                       |From new raw data                                                                                                                                                  
 210   |22.5 GHz (VLA)      |2.1E+01               |+/-1         |milliJy             |2.25E+10 |2.10E-02    |1.0E-03                   |1.0E-03                   |                           |                           |+/-1.00E-03    |Jy       |2008A&A...477...95C|uncertainty            |22.5 GHz           |Broad-band measurement                                                 |04 34 00.02 -08 34 44.98 (J2000)|Flux integrated from map                                |                                       |From new raw data                                                                                                                                                  
 211   |10.63 GHz (ARO)     |3.0E+01               |+/-13        |milliJy             |1.06E+10 |3.00E-02    |1.3E-02                   |1.3E-02                   |                           |                           |+/-1.30E-02    |Jy       |1995ApJS...98..369B|rms uncertainty        |10.63 GHz          |Broad-band measurement                                                 |                                |Flux integrated from map                                |Probable detection                     |From new raw data                                                                                                                                                  
 212   |8.46 GHz (VLA)      |4.1E+01               |+/-0.6       |milliJy             |8.46E+09 |4.11E-02    |6.0E-04                   |6.0E-04                   |                           |                           |+/-6.00E-04    |Jy       |2006ApJS..164...52S|uncertainty            |8.46   GHz         |Broad-band measurement                                                 |04 34 00.0 -08 34 45 (J2000)    |Flux integrated from map                                |                                       |From new raw data                                                                                                                                                  
 213   |4.85 GHz            |6.3E+01               |+/-11        |milliJy             |4.85E+09 |6.30E-02    |1.1E-02                   |1.1E-02                   |                           |                           |+/-1.10E-02    |Jy       |1995ApJS...97..347G|rms noise              |4.85       GHz     |Broad-band measurement                                                 |043402.5 -083444 (J2000)        |Modelled datum                                          |                                       |From new raw data; Corrected for contaminating sources                                                                                                             
 214   |4.755 GHz (GBT)     |6.4E+01               |+/-6         |milliJy             |4.76E+09 |6.40E-02    |6.0E-03                   |6.0E-03                   |                           |                           |+/-6.00E-03    |Jy       |1995ApJS...98..369B|rms uncertainty        |4.755 GHz          |Broad-band measurement                                                 |                                |Flux integrated from map                                |Probable detection                     |From new raw data                                                                                                                                                  
 217   |1398 MHz (VLA)      |1.4E+02               |             |milliJy             |1.40E+09 |1.40E-01    |                          |                          |                           |                           |               |Jy       |2010A&A...513A..11O|no uncertainty reported|1398 GHz           |Broad-band measurement                                                 |04 34 00.06 -08 34 44.6 (J2000) |Total flux                                              |Flux in central region                 |From new raw data                                                                                                                                                  
 218   |1.4GHz              |1.4E+02               |+/-4.9       |milliJy             |1.40E+09 |1.38E-01    |4.9E-03                   |4.9E-03                   |                           |                           |+/-4.90E-03    |Jy       |1998AJ....115.1693C|uncertainty            |1.40   GHz         |Broad-band measurement                                                 |04 34 0.02 -08 34 45.1 (J2000)  |Flux integrated from map                                |                                       |From new raw data                                                                                                                                                  
 219   |610 MHz (GMRT)      |2.0E-01               |+/-0.005     |Jy                  |6.10E+08 |2.02E-01    |5.0E-03                   |5.0E-03                   |                           |                           |+/-5.00E-03    |Jy       |2010MNRAS.405..887C|uncertainty            |610 MHz            |Broad-band measurement                                                 |                                |Flux integrated from map                                |                                       |From new raw data                                                                                                                                                  
 220   |244 MHz (GMRT)      |2.5E-01               |+/-0.040     |Jy                  |2.44E+08 |2.50E-01    |4.0E-02                   |4.0E-02                   |                           |                           |+/-4.00E-02    |Jy       |2010MNRAS.405..887C|uncertainty            |244 MHz            |Broad-band measurement                                                 |                                |Flux integrated from map                                |                                       |From new raw data                                                                                                                                                  
