
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2016-06-16T17:03:17PDT



Photometric Data for PKS 1623+26:[SSP2004] BX0663

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|G (WHT)             | 24.38     ||mag                 |6.38E+14|  6.43E-07||Jy|2006ApJ...647..128E|no uncertainty reported|    0.47   microns   | Broad-band measurement|| Flux in fixed aperture|                                        |Averaged from previously published data
2|H{alpha} (Keck II)  | 8.2E-17   |+/-0.3E-17|erg s^-1^ cm^-2^    |4.57E+14|  8.20E+06|+/-3.00E+05|Jy-Hz|2006ApJ...646..107E|uncertainty|    6563   A         | Line measurement; flux integrated over line; lines measured in emission|16 26 04.58 +26 48 00.20 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
3|H{alpha} (Keck)     | 16.8E-17  |+/-0.9E-17| erg/s/cm^2^        |4.57E+14|  1.68E+07|+/-9.00E+05|Jy-Hz|2004ApJ...612..108S|internal error|      6563 A         | Line measurement; flux integrated over line; lines measured in emission|16 26 04.576 26 48 00.202 (J2000)| Flux integrated from map|Double-peaked emission line             |From new raw data
4|H{alpha} (VLT)      | 16.7E-17  |+/-0.9E-17|erg/s/cm^2^         |4.57E+14|  1.67E+07|+/-9.00E+05|Jy-Hz|2009ApJ...706.1364F|uncertainty|      6563 A         | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|                                        |From new raw data
5|[N II] (Keck)       | 3.5E-17   |+/-0.3E-17| erg/s/cm^2^        |4.55E+14|  3.50E+06|+/-3.00E+05|Jy-Hz|2004ApJ...612..108S|internal error|      6584 A         | Line measurement; flux integrated over line; lines measured in emission|16 26 04.576 26 48 00.202 (J2000)| Flux integrated from map|                                        |From new raw data
6|J (Hale/WIRC)       | 22.51     ||mag                 |2.40E+14|  1.55E-06||Jy|2006ApJ...646..107E|no uncertainty reported|    1.25   microns   | Broad-band measurement|16 26 04.58 +26 48 00.20 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data; derived from aflux in a different band and a color
7|F160W (HST) AB      | 22.79     |+/-0.10 |mag                 |1.87E+14|  2.78E-06|+/-2.56E-07|Jy|2011ApJ...731...65F|uncertainty|     1.603 microns   | Broad-band measurement|| Flux in fixed aperture|                                        |From new raw data
8|K_s (Hale/WIRC)     | 19.92     ||mag                 |1.39E+14|  7.21E-06||Jy|2006ApJ...646..107E|no uncertainty reported|    2.15   microns   | Broad-band measurement|16 26 04.58 +26 48 00.20 (J2000)| Flux in fixed aperture|                                        |Averaged new and previously published data
9|CO(3-2) (PdBI)      |           |+/-0.18 |Jy km/s             |3.46E+11||+/-6.06E+04|Jy-Hz|2010Natur.463..781T|1 sigma|   345.998 GHz       | Line measurement; flux integrated over line; lines measured in emission|| Flux integrated from map|                                        |From new raw data
