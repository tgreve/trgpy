
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-05-27T08:07:49PDT



Photometric Data for GN 850.07

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|2-8 keV (Chandra)   | |<17.4E-17  |erg/cm^2^/s         |1.21E+18| |1.44E-11|Jy|2009ApJ...698.1380M|no uncertainty reported|      5.00 keV       | Broad-band measurement|12 36 21.27 +62 17 08.1 (J2000)| Not reported in paper|                                        |Averaged from previously published data; NED frequencyassigned to mid-point of band in keV
2|0.5-8 keV (Chandra) | |<10.9E-17  |erg/cm^2^/s         |1.03E+18| |1.06E-11|Jy|2009ApJ...698.1380M|no uncertainty reported|      4.25 keV       | Broad-band measurement|12 36 21.27 +62 17 08.1 (J2000)| Not reported in paper|                                        |Averaged from previously published data; NED frequencyassigned to mid-point of band in keV
3|H{alpha} (Keck)     | 2.0E-19   |+/-0.6E-19| W/m^2^             |4.57E+14|  2.00E+07|+/-6.00E+06|Jy-Hz|2004ApJ...617...64S|uncertainty|      6563 A         | Line measurement; flux integrated over line; lines measured in emission|123621.27 +621708.4 (J2000)| Flux integrated from map|                                        |From new raw data
4|I (Cousins)         | 24.92     |+/-0.15 |mag                 |3.79E+14|  2.75E-07|+/-4.07E-08|Jy|2004ApJ...616...71S|1 sigma|    7900   A         | Broad-band measurement| | Flux in fixed aperture|4" aper; phot contam by near neighbor   |Averaged new and previously published data
6|K_s (Hale/WIRC) AB  | 22.44     | |mag                 |1.39E+14|  3.84E-06| |Jy|2005ApJ...633..748R|no uncertainty reported|   2.150   microns   | Broad-band measurement|12 36 21.27 +62 17 08.4 (J2000)| Flux in fixed aperture|                                        |From new raw data
7|K_s_ (2MASS)        | 20.73     |+/-0.33 |mag                 |1.38E+14|  3.40E-06|+/-1.21E-06|Jy|2004ApJ...616...71S|1 sigma|    2.17   microns   | Broad-band measurement| | Flux in fixed aperture|4" aper; phot contam by near neighbor   |Averaged new and previously published data
8|3.6 microns (IRAC)  | 13.3      |+/-1.6  |microJy             |8.44E+13|  1.33E-05|+/-1.60E-06|Jy|2009ApJ...699.1610H|uncertainty|     3.550 microns   | Broad-band measurement|12 36 21.34 +62 17 08.3 (J2000)| Flux in fixed aperture|                                        |From new raw data
9|4.5 microns (IRAC)  | 20.0      |+/-2.2  |microJy             |6.67E+13|  2.00E-05|+/-2.20E-06|Jy|2009ApJ...699.1610H|uncertainty|     4.493 microns   | Broad-band measurement|12 36 21.34 +62 17 08.3 (J2000)| Flux in fixed aperture|                                        |From new raw data
10|5.8 microns (IRAC)  | 23.5      |+/-3.4  |microJy             |5.23E+13|  2.35E-05|+/-3.40E-06|Jy|2009ApJ...699.1610H|uncertainty|     5.731 microns   | Broad-band measurement|12 36 21.34 +62 17 08.3 (J2000)| Flux in fixed aperture|                                        |From new raw data
11|8.0 microns (IRAC)  | 19.3      |+/-2.1  |microJy             |3.85E+13|  1.93E-05|+/-2.10E-06|Jy|2009ApJ...699.1610H|uncertainty|     7.782 microns   | Broad-band measurement|12 36 21.34 +62 17 08.3 (J2000)| Flux in fixed aperture|                                        |From new raw data
12|16 microns (Spitzer)| |<30.0      |microJy             |1.87E+13| |3.00E-05|Jy|2009ApJ...698.1380M|no uncertainty reported|        16 microns   | Broad-band measurement|12 36 21.27 +62 17 08.1 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
13|16 microns (Spitzer)| 0.048     |+/-0.007| milliJy            |1.87E+13|  4.80E-05|+/-7.00E-06|Jy|2008ApJ...675.1171P|uncertainty|        16 microns   | Broad-band measurement|12 36 21.27 +62 17 08.1 (J2000)| Flux integrated from map|                                        |Averaged from previously published data
14|24 microns (IRAC)   | 370.0     |+/-11.4 | microJy            |1.27E+13|  3.70E-04|+/-1.14E-05|Jy|2009ApJ...691..560C|uncertainty|     23.68 microns   | Broad-band measurement|12 36 21.25 +62 17 08.3 (J2000)| Not reported in paper|                                        |Averaged from previously published data
15|24 microns (Spitzer)| 347       | |microJy             |1.27E+13|  3.47E-04| |Jy|2009ApJ...698.1380M|no uncertainty reported|     23.68 microns   | Broad-band measurement|12 36 21.27 +62 17 08.1 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
16|24 microns (MIPS)   | 357.0     |+/-38.0 |microJy             |1.27E+13|  3.57E-04|+/-3.80E-05|Jy|2009ApJ...699.1610H|uncertainty|     23.68 microns   | Broad-band measurement|123621.27 +621708.4 (J2000)| Flux in fixed aperture|                                        |From new raw data
17|70 microns (Spitzer)| |<3.5       | milliJy            |4.20E+12| |3.50E-03|Jy|2008ApJ...675.1171P|3rms uncertainty reported|     71.42 microns   | Broad-band measurement|12 36 21.27 +62 17 08.1 (J2000)| Flux integrated from map|                                        |Averaged from previously published data
18|70 microns (Spitzer)| |<3000      |microJy             |4.20E+12| |3.00E-03|Jy|2009ApJ...698.1380M|3rms uncertainty reported|     71.42 microns   | Broad-band measurement|12 36 21.27 +62 17 08.1 (J2000)| Flux in fixed aperture|                                        |Averaged from previously published data
19|70 microns (MIPS)   | |<2.2       |microJy             |4.20E+12| |2.20E-03|Jy|2009ApJ...699.1610H|3 sigma|     71.42 microns   | Broad-band measurement|123621.27 +621708.4 (J2000)| Flux in fixed aperture|                                        |From new raw data
20|850 microns (SCUBA) | 8.9       |+/-1.5  |milliJy             |3.53E+11|  8.90E-03|+/-1.50E-03|Jy|2005MNRAS.358..149P|uncertainty|     850   microns   | Broad-band measurement|12 36 21.3 +62 17 11 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
21|850 microns (SCUBA) | 7.8       |+/-1.9  |milliJy             |3.53E+11|  7.80E-03|+/-1.90E-03|Jy|2005ApJ...622..772C|uncertainty|     850   microns   | Broad-band measurement|123621.27 +621708.4 (J2000)| Flux integrated from map|                                        |From new raw data
22|1.4 GHz (VLA)       | 138       |+/-7    | microJy            |1.40E+09|  1.38E-04|+/-7.00E-06|Jy|2006MNRAS.371..963B|1 sigma|       1.4 GHz       | Broad-band measurement|12 36 21.272 +62 17 08.36 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
23|1.4 GHz (VLA)       | 169.4     |+/-8.8  | microJy            |1.40E+09|  1.69E-04|+/-8.80E-06|Jy|2009ApJ...691..560C|uncertainty|       1.4 GHz       | Broad-band measurement|12 36 21.25 +62 17 08.3 (J2000)| Not reported in paper|                                        |From reprocessed raw data
24|1.4 GHz             | 148.0     |+/-11.0 |microJy             |1.40E+09|  1.48E-04|+/-1.10E-05|Jy|2000ApJ...533..611R|1 sigma|1.4        GHz       | Broad-band measurement; broad-band flux derived by integration over spectrum; synthetic band|123621.272 +621708.40 (J2000)| Flux integrated from map; Pointing and beam filling|                                        |From new raw data; Corrected for contaminating sources
25|1.4 GHz (VLA)       | 148       | |microJy             |1.40E+09|  1.48E-04| |Jy|2005MNRAS.358.1159M|no uncertainty reported|     1.4   GHz       | Broad-band measurement|12 36 21.2691 +62 17 08.458 (J2000)| Flux integrated from map|                                        |From new raw data
26|1.4 GHz (VLA)       | 162.9     |+/-7.0  |microJy             |1.40E+09|  1.63E-04|+/-7.00E-06|Jy|2010ApJS..188..178M|uncertainty|       1.4 GHz       | Broad-band measurement|12 36 21.25 +62 17 08.3 (J2000)| Total flux; Beam filling or dilution corrected|Major=0.0"; Minor=0.0"; PA=0 deg        |From new raw data
