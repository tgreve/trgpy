\queryDateTime = 2018-11-26T07:47:29PST
\source = /hydra/workarea/irsaviewer/temp_files/IpacTableFromSource2927304954651768398.tbl
\QUERY_STATUS = OK
\CatalogTargetColName = Coordinates Targeted
\Description = Published and Homogenized [Frequency, Flux Dens...
\LINK = http://ned.ipac.caltech.edu/cgi-bin/datasearch?sea
\
z=0.00379
|No.   |Observed Passband   |Photometry Measurement|Uncertainty  |Units               |Frequency|Flux Density|Upper limit of uncertainty|Lower limit of uncertainty|Upper limit of Flux Density|Lower limit of Flux Density|NED Uncertainty|NED Units|Refcode            |Significance                  |Published frequency|Frequency Mode                                                         |Coordinates Targeted             |Spatial Mode                                            |Qualifiers                              |Comments                                                                                                                                                           |
|int   |char                |double                |char         |char                |double   |double      |double                    |double                    |double                     |double                     |char           |char     |char               |char                          |char               |char                                                                   |char                             |char                                                    |char                                    |char                                                                                                                                                               |
|      |                    |                      |             |                    |Hz       |Jy          |                          |                          |                           |                           |               |         |                   |                              |                   |                                                                       |                                 |                                                        |                                        |                                                                                                                                                                   |
|      |                    |                      |             |                    |         |            |                          |                          |                           |                           |               |         |                   |                              |                   |                                                                       |                                 |                                                        |                                        |                                                                                                                                                                   |
 1     |0.1-100 GeV (Fermi) |5.7E-12               |+/-1.2E-12   |erg/cm^2^/s         |1.21E+25 |4.71E-14    |9.92E-15                  |9.92E-15                  |                           |                           |+/-9.92E-15    |Jy       |2012ApJS..199...31N|1 sigma                       |50.05 GeV          |Broad-band measurement                                                 |040.650 +00.104 (J2000)          |Modelled datum                                          |                                        |From new raw data; NED frequency assigned to mid-point ofband in keV                                                                                               
 2     |14-195 keV (Swift)  |3.7E-11               |+/-0.53E-11  |erg/s/cm^2^         |2.53E+19 |1.47E-07    |2.09E-08                  |2.09E-08                  |                           |                           |+/-2.09E-08    |Jy       |2010ApJS..186..378T|uncertainty                   |104.50 keV         |Broad-band measurement                                                 |040.638 +00.000 (J2000)          |Flux integrated from map                                |                                        |From new raw data; NED frequency assigned to mid-point ofband in keV                                                                                               
 3     |15-150 keV (Swift)  |2.7E-11               |+/-5.4e-12   |erg/cm^2^/s         |1.99E+19 |1.36E-07    |2.71E-08                  |2.71E-08                  |                           |                           |+/-2.71E-08    |Jy       |2010A&A...524A..64C|uncertainty                   |82.50 keV          |Broad-band measurement                                                 |040.671 -00.017 (J2000)          |Modelled datum                                          |                                        |From new raw data; NED frequency assigned to mid-point ofband in keV                                                                                               
 4     |40-100 keV INTEGRAL |1.7E-11               |+/-0.48E-11  |erg cm^-2^ s^-1^    |1.69E+19 |9.82E-08    |2.84E-08                  |2.84E-08                  |                           |                           |+/-2.84E-08    |Jy       |2006ApJ...638..642B|uncertainty                   |70   keV           |Broad-band measurement                                                 |02 42 41 -00 00 48 (J2000)       |Flux integrated from map                                |                                        |From new raw data; NED frequency assigned to mid-point ofband in keV                                                                                               
 5     |40-100 keV INTEGRAL |1.9E+00               |+/-0.4       |milliCrab           |1.69E+19 |1.06E-07    |2.23E-08                  |2.23E-08                  |                           |                           |+/-2.23E-08    |Jy       |2007ApJS..170..175B|uncertainty                   |70   keV           |Broad-band measurement                                                 |040.689 +00.016 (J2000)          |Flux integrated from map                                |Time-averaged flux                      |From reprocessed raw data; NED frequency assigned tomid-point of band in keV                                                                                       
 6     |40-100 keV INTEGRAL |1.3E-11               |             |erg/cm^2^/s         |1.69E+19 |7.51E-08    |                          |                          |                           |                           |               |Jy       |2009A&A...505..417B|no uncertainty reported       |70.00 keV          |Broad-band measurement                                                 |40.67012 -0.01344 (J2000)        |Modelled datum                                          |                                        |From new raw data; NED frequency assigned to mid-point ofband in keV                                                                                               
 7     |20-100 keV INTEGRAL |3.0E-11               |             |erg/s/cm^2^         |1.45E+19 |2.07E-07    |                          |                          |                           |                           |               |Jy       |2009MNRAS.399..944M|no uncertainty reported       |60.00 keV          |Broad-band measurement                                                 |02 42 40.71 -00 00 47.8 (J2000)  |Flux integrated from map                                |                                        |Averaged from previously published data; NED frequencyassigned to mid-point of band in keV                                                                         
 8     |17-80 keV (INTEGRAL)|1.9E-11               |+/-1.23E-11  |erg/cm^2^/s         |1.17E+19 |1.59E-07    |1.05E-07                  |1.05E-07                  |                           |                           |+/-1.05E-07    |Jy       |2010A&A...524A..72L|uncertainty                   |48.5  keV          |Broad-band measurement                                                 |                                 |Modelled datum                                          |                                        |From new raw data; NED frequency assigned to mid-point ofband in keV                                                                                               
 9     |17-60 keV (INTEGRAL)|1.9E-11               |+/-0.30E-11  |erg s^-1^ cm^-2^    |9.31E+18 |2.04E-07    |3.22E-08                  |3.22E-08                  |                           |                           |+/-3.22E-08    |Jy       |2007A&A...462...57S|uncertainty                   |38.50   keV        |Broad-band measurement                                                 |                                 |Flux integrated from map                                |                                        |Averaged new and previously published data; NED frequencyassigned to mid-point of band in keV                                                                      
 10    |15-55 keV (Swift)   |2.0E-11               |+/-0.22E-11  |erg/cm^2^/s         |8.46E+18 |2.36E-07    |2.60E-08                  |2.60E-08                  |                           |                           |+/-2.60E-08    |Jy       |2009ApJ...699..603A|uncertainty                   |35.00 keV          |Broad-band measurement                                                 |040.732 -00.012 (J2000)          |Flux integrated from map                                |                                        |From reprocessed raw data; NED frequency assigned tomid-point of band in keV                                                                                       
 11    |20-40 keV (INTEGRAL)|9.3E-12               |+/-0.27E-11  |erg cm^-2^ s^-1^    |7.25E+18 |1.28E-07    |3.72E-08                  |3.72E-08                  |                           |                           |+/-3.72E-08    |Jy       |2006ApJ...638..642B|uncertainty                   |30   keV           |Broad-band measurement                                                 |02 42 41 -00 00 48 (J2000)       |Flux integrated from map                                |                                        |From new raw data; NED frequency assigned to mid-point ofband in keV                                                                                               
 12    |20-40 keV (INTEGRAL)|1.6E+00               |+/-0.2       |milliCrab           |7.25E+18 |1.67E-07    |2.09E-08                  |2.09E-08                  |                           |                           |+/-2.09E-08    |Jy       |2007ApJS..170..175B|uncertainty                   |30   keV           |Broad-band measurement                                                 |040.689 +00.016 (J2000)          |Flux integrated from map                                |Time-averaged flux                      |From reprocessed raw data; NED frequency assigned tomid-point of band in keV                                                                                       
 13    |20-40 keV (INTEGRAL)|1.2E-11               |             |erg/cm^2^/s         |7.25E+18 |1.60E-07    |                          |                          |                           |                           |               |Jy       |2009A&A...505..417B|no uncertainty reported       |30.00 keV          |Broad-band measurement                                                 |40.67012 -0.01344 (J2000)        |Modelled datum                                          |                                        |From new raw data; NED frequency assigned to mid-point ofband in keV                                                                                               
 14    |10-50 keV (Suzaku)  |1.4E+00               |             |log(erg/s/cm^2^)    |7.25E+18 |3.39E-07    |                          |                          |                           |                           |               |Jy       |2011ApJ...727...19F|no uncertainty reported       |30.00 keV          |Broad-band measurement                                                 |                                 |Modelled datum                                          |                                        |From reprocessed raw data; NED frequency assigned tomid-point of band in keV                                                                                       
 15    |3.5-15 keV (XMM)    |6.3E-12               |             |erg cm^-2^ s^-1^    |2.24E+18 |2.81E-07    |                          |                          |                           |                           |               |Jy       |2006MNRAS.368..707P|no uncertainty reported       |9.25   keV         |Broad-band measurement                                                 |                                 |Flux integrated from map                                |                                        |From new raw data; NED frequency assigned to mid-point ofband in keV                                                                                               
 16    |F_2-10_ keV         |5.3E-01               |+/-10  %     |10^-11^ erg/s/cm^2^ |1.45E+18 |3.65E-07    |3.65E-08                  |3.65E-08                  |                           |                           |+/-3.65E-08    |Jy       |1989MNRAS.240..833T|typical accuracy              |6.0    keV         |Broad-band measurement                                                 |                                 |Flux integrated from map                                |Energy index 0.72                       |From new raw data; NED frequency assigned to mid-point ofband in keV                                                                                               
 17    |2-10 keV (XMM)      |4.6E-12               |             |erg cm^-2^ s^-1^    |1.45E+18 |3.19E-07    |                          |                          |                           |                           |               |Jy       |2006A&A...446..459C|no uncertainty reported       |6   keV            |Broad-band measurement                                                 |02 42 40.7 -00 00 47.6 (J2000)   |Flux integrated from map                                |                                        |From new raw data; Uncorrected for known sources in beam; NEDfrequency assigned to mid-point of band in keV                                                        
 18    |2-10 keV            |3.5E-15               |             |W/m^2^              |1.45E+18 |2.41E-07    |                          |                          |                           |                           |               |Jy       |2004A&A...418..465L|no uncertainty reported       |6   keV            |Broad-band measurement                                                 |                                 |Flux integrated from map                                |Observed flux                           |Averaged from previously published data; NED frequencyassigned to mid-point of band in keV                                                                         
 19    |2-10 keV (ASCA)     |3.7E-12               |             |ergs/s/cm^2^        |1.45E+18 |2.58E-07    |                          |                          |                           |                           |               |Jy       |2001ApJS..133....1U|no uncertainty reported       |6.00 keV           |Broad-band measurement                                                 |040.6719 -00.0054 (J2000)        |Flux integrated from map                                |                                        |From reprocessed raw data; Extinction-corrected for MilkyWay; NED frequency assigned to mid-point of band in keV                                                   
 20    |2-10 keV            |5.4E-12               |+/-110E-13   |erg/s/cm^2^         |1.45E+18 |3.74E-07    |7.59E-07                  |7.59E-07                  |                           |                           |+/-7.59E-07    |Jy       |2011ApJ...729...52L|uncertainty                   |6.00 keV           |Broad-band measurement                                                 |                                 |Modelled datum                                          |                                        |From reprocessed raw data; NED frequency assigned tomid-point of band in keV                                                                                       
 21    |2-10 keV (Chandra)  |5.6E-12               |             |erg/cm^2^/s         |1.45E+18 |3.86E-07    |                          |                          |                           |                           |               |Jy       |2011ApJ...738..147S|no uncertainty reported       |6.00 keV           |Broad-band measurement                                                 |                                 |Modelled datum                                          |                                        |From reprocessed raw data; NED frequency assigned tomid-point of band in keV                                                                                       
 22    |2-10 keV (XMM)      |5.0E-12               |             |erg/s/cm^2^         |1.45E+18 |3.43E-07    |                          |                          |                           |                           |               |Jy       |2011MNRAS.413.1206B|no uncertainty reported       |6.00 keV           |Broad-band measurement                                                 |040.672 -00.013 (J2000)          |Modelled datum                                          |                                        |From reprocessed raw data; NED frequency assigned tomid-point of band in keV                                                                                       
 23    |2-8 keV (ASCA)      |5.2E-12               |             |ergs/cm^2^/s        |1.21E+18 |4.29E-07    |                          |                          |                           |                           |               |Jy       |2007AJ....134.1263C|no uncertainty reported       |5.00 keV           |Broad-band measurement                                                 |                                 |Modelled datum                                          |                                        |Averaged from previously published data; NED frequencyassigned to mid-point of band in keV                                                                         
 24    |0.3-8 keV (Chandra) |1.8E-11               |             |erg/s/cm^2^         |1.00E+18 |1.79E-06    |                          |                          |                           |                           |               |Jy       |2011ApJS..192...10L|no uncertainty reported       |4.15 keV           |Broad-band measurement                                                 |02 42 40.793 -00 00 46.44 (J2000)|Flux integrated from map                                |                                        |From reprocessed raw data; NED frequency assigned tomid-point of band in keV                                                                                       
 25    |0.7-7 keV (ASCA)    |8.8E-12               |             |ergs/s/cm^2^        |9.31E+17 |9.47E-07    |                          |                          |                           |                           |               |Jy       |2001ApJS..133....1U|no uncertainty reported       |3.85 keV           |Broad-band measurement                                                 |040.6719 -00.0054 (J2000)        |Flux integrated from map                                |                                        |From reprocessed raw data; Extinction-corrected for MilkyWay; NED frequency assigned to mid-point of band in keV                                                   
 26    |0.2-4 keV (EINSTEIN)|2.1E-11               |             |ergs sec^-1^ cm^-2^ |5.25E+17 |3.94E-06    |                          |                          |                           |                           |               |Jy       |1992ApJS...80..531F|no uncertainty reported       |2.1    keV         |Broad-band measurement; synthetic band                                 |02 40 07 -00 13 27 (B1950)       |Flux integrated from map                                |                                        |From reprocessed raw data; Extinction-corrected for MilkyWay; NED frequency assigned to mid-point of band in keV                                                   
 27    |0.3-3 keV (XMM)     |1.6E-11               |             |erg cm^-2^ s^-1^    |3.99E+17 |4.01E-06    |                          |                          |                           |                           |               |Jy       |2006MNRAS.368..707P|no uncertainty reported       |1.65   keV         |Broad-band measurement                                                 |                                 |Flux integrated from map                                |                                        |From new raw data; NED frequency assigned to mid-point ofband in keV                                                                                               
 28    |0.7-2 keV (ASCA)    |5.8E-12               |             |ergs/s/cm^2^        |3.26E+17 |1.78E-06    |                          |                          |                           |                           |               |Jy       |2001ApJS..133....1U|no uncertainty reported       |1.35 keV           |Broad-band measurement                                                 |040.6719 -00.0054 (J2000)        |Flux integrated from map                                |                                        |From reprocessed raw data; Extinction-corrected for MilkyWay; NED frequency assigned to mid-point of band in keV                                                   
 29    |0.1-2.4 keV (ROSAT) |3.6E-11               |+/-1.66E-12  |ergs sec^-1^ cm^-2^ |3.25E+17 |1.09E-05    |5.11E-07                  |5.11E-07                  |                           |                           |+/-5.11E-07    |Jy       |1994A&A...281..355B|based on count statistics only|1.3   keV          |Broad-band measurement; synthetic band                                 |                                 |Flux integrated from map                                |                                        |From new raw data; Extinction-corrected for Milky Way                                                                                                              
 30    |0.5-2 keV (XMM)     |1.1E-11               |             |erg cm^-2^ s^-1^    |3.02E+17 |3.69E-06    |                          |                          |                           |                           |               |Jy       |2006A&A...446..459C|no uncertainty reported       |1.25   keV         |Broad-band measurement                                                 |02 42 40.7 -00 00 47.6 (J2000)   |Flux integrated from map                                |                                        |From new raw data; Uncorrected for known sources in beam; NEDfrequency assigned to mid-point of band in keV                                                        
 31    |0.5-2 keV (ASCA)    |1.0E-11               |             |ergs/cm^2^/s        |3.02E+17 |3.38E-06    |                          |                          |                           |                           |               |Jy       |2007AJ....134.1263C|no uncertainty reported       |1.25 keV           |Broad-band measurement                                                 |                                 |Modelled datum                                          |                                        |Averaged from previously published data; NED frequencyassigned to mid-point of band in keV                                                                         
 33    |1030 A (FUSE)       |2.3E-14               |             |erg/cm^2^/s/A       |2.91E+15 |8.15E-04    |                          |                          |                           |                           |               |Jy       |2006ApJS..165..229F|no uncertainty reported       |1030   A           |Broad-band measurement                                                 |                                 |Flux integrated from map                                |S/N = 29.3                              |From reprocessed raw data                                                                                                                                          
 34    |1482A (IUE)         |6.6E-14               |+/-1.06E-14  |ergs cm^-2 s^-1 A^-1|2.02E+15 |4.87E-03    |7.78E-04                  |7.78E-04                  |                           |                           |+/-7.78E-04    |Jy       |1993ApJS...86....5K|uncertainty                   |1482   A           |Broad-band measurement; flux integrated over line                      |                                 |Flux in fixed aperture                                  |20"x10" aperture                        |Averaged from new and transformed previously published data                                                                                                        
 35    |FUV (GALEX) AB      |1.3E+01               |+/-0.01      |mag                 |1.98E+15 |2.78E-02    |2.56E-04                  |2.56E-04                  |                           |                           |+/-2.56E-04    |Jy       |2007ApJS..173..185G|uncertainty                   |1516 A             |Broad-band measurement                                                 |02 42 40.7 -00 00 47.8 (J2000)   |Total flux                                              |                                        |From new raw data                                                                                                                                                  
 36    |FUV (GALEX) AB      |1.5E+01               |             |mag                 |1.98E+15 |3.10E-03    |                          |                          |                           |                           |               |Jy       |2007ApJS..173..404B|no uncertainty reported       |1516 A             |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |                                        |From reprocessed raw data; Extinction-corrected for Milky Way                                                                                                      
 37    |FUV (GALEX) AB      |1.3E+01               |+/-0.10      |mag                 |1.96E+15 |3.33E-02    |3.06E-03                  |3.06E-03                  |                           |                           |+/-3.06E-03    |Jy       |2014ApJS..212...18B|uncertainty                   |1531   A           |Broad-band measurement                                                 |40.66969000 -0.01318000 (J2000)  |Flux in fixed aperture                                  |155"x180" aperture                      |From new raw data; Extinction-corrected for Milky Way                                                                                                              
 38    |FUV (GALEX) AB      |1.3E+01               |+/-0.10      |mag                 |1.96E+15 |2.30E-02    |2.12E-03                  |2.12E-03                  |                           |                           |+/-2.12E-03    |Jy       |2014ApJS..212...18B|uncertainty                   |1531   A           |Broad-band measurement                                                 |40.66969000 -0.01318000 (J2000)  |Flux in fixed aperture                                  |155"x180" aperture                      |From new raw data                                                                                                                                                  
 39    |1550 A (OAO)        |1.0E+01               |+/-0.64      |mag                 |1.93E+15 |2.42E-02    |1.95E-02                  |1.95E-02                  |                           |                           |+/-1.95E-02    |Jy       |1982ApJ...256....1C|rms noise                     |1550       A       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |Aperture 10.0 arcmin                    |From new raw data                                                                                                                                                  
 40    |1910 A (OAO)        |1.0E+01               |+/-0.78      |mag                 |1.57E+15 |3.06E-02    |3.22E-02                  |3.22E-02                  |                           |                           |+/-3.22E-02    |Jy       |1982ApJ...256....1C|rms noise                     |1910       A       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |Aperture 10.0 arcmin                    |From new raw data                                                                                                                                                  
 41    |1913A (IUE)         |7.5E-14               |+/-3.00E-14  |ergs cm^-2 s^-1 A^-1|1.57E+15 |9.20E-03    |3.67E-03                  |3.67E-03                  |                           |                           |+/-3.67E-03    |Jy       |1993ApJS...86....5K|uncertainty                   |1913   A           |Broad-band measurement; flux integrated over line                      |                                 |Flux in fixed aperture                                  |20"x10" aperture                        |Averaged from new and transformed previously published data                                                                                                        
 42    |NUV (GALEX) AB      |1.2E+01               |+/-0.01      |mag                 |1.32E+15 |4.70E-02    |4.33E-04                  |4.33E-04                  |                           |                           |+/-4.33E-04    |Jy       |2007ApJS..173..185G|uncertainty                   |2267 A             |Broad-band measurement                                                 |02 42 40.7 -00 00 47.8 (J2000)   |Total flux                                              |                                        |From new raw data                                                                                                                                                  
 43    |NUV (GALEX) AB      |1.2E+01               |+/-0.10      |mag                 |1.31E+15 |4.39E-02    |4.05E-03                  |4.05E-03                  |                           |                           |+/-4.05E-03    |Jy       |2014ApJS..212...18B|uncertainty                   |2286   A           |Broad-band measurement                                                 |40.66969000 -0.01318000 (J2000)  |Flux in fixed aperture                                  |155"x180" aperture                      |From new raw data                                                                                                                                                  
 44    |NUV (GALEX) AB      |1.2E+01               |+/-0.10      |mag                 |1.31E+15 |6.38E-02    |5.88E-03                  |5.88E-03                  |                           |                           |+/-5.88E-03    |Jy       |2014ApJS..212...18B|uncertainty                   |2286   A           |Broad-band measurement                                                 |40.66969000 -0.01318000 (J2000)  |Flux in fixed aperture                                  |155"x180" aperture                      |From new raw data; Extinction-corrected for Milky Way                                                                                                              
 45    |2373A (IUE)         |5.5E-14               |+/-1.54E-14  |ergs cm^-2 s^-1 A^-1|1.26E+15 |1.04E-02    |2.90E-03                  |2.90E-03                  |                           |                           |+/-2.90E-03    |Jy       |1993ApJS...86....5K|uncertainty                   |2373   A           |Broad-band measurement; flux integrated over line                      |                                 |Flux in fixed aperture                                  |20"x10" aperture                        |Averaged from new and transformed previously published data                                                                                                        
 46    |2460 A (OAO)        |1.1E+01               |+/-0.54      |mag                 |1.22E+15 |4.03E-02    |2.60E-02                  |2.60E-02                  |                           |                           |+/-2.60E-02    |Jy       |1982ApJ...256....1C|rms noise                     |2460       A       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |Aperture 10.0 arcmin                    |From new raw data                                                                                                                                                  
 47    |2700A (IUE)         |4.8E-14               |+/-0.20E-14  |ergs cm^-2 s^-1 A^-1|1.11E+15 |1.17E-02    |4.87E-04                  |4.87E-04                  |                           |                           |+/-4.87E-04    |Jy       |1993ApJS...86....5K|uncertainty                   |2700   A           |Broad-band measurement; flux integrated over line                      |                                 |Flux in fixed aperture                                  |20"x10" aperture                        |Averaged from new and transformed previously published data                                                                                                        
 48    |2980 A (OAO)        |1.0E+01               |+/-0.13      |mag                 |1.01E+15 |1.10E-01    |1.40E-02                  |1.40E-02                  |                           |                           |+/-1.40E-02    |Jy       |1982ApJ...256....1C|rms noise                     |2980       A       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |Aperture 10.0 arcmin                    |From new raw data                                                                                                                                                  
 49    |3320 A (OAO)        |9.7E+00               |+/-0.03      |mag                 |9.03E+14 |1.78E-01    |4.98E-03                  |4.98E-03                  |                           |                           |+/-4.98E-03    |Jy       |1982ApJ...256....1C|rms noise                     |3320       A       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |Aperture 10.0 arcmin                    |From new raw data                                                                                                                                                  
 50    |3390A               |1.2E+00               |+/-10  %     |10^-26 erg/cm^2/s/Hz|8.85E+14 |1.21E-02    |1.21E-03                  |1.21E-03                  |                           |                           |+/-1.21E-03    |Jy       |1970ApJ...162..743A|estimated error               |3390       A       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |8" aperture                             |From new raw data                                                                                                                                                  
 51    |3448A               |1.5E+00               |+/-10  %     |10^-26 erg/cm^2/s/Hz|8.70E+14 |1.54E-02    |1.54E-03                  |1.54E-03                  |                           |                           |+/-1.54E-03    |Jy       |1970ApJ...162..743A|estimated error               |3448       A       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |8" aperture                             |From new raw data                                                                                                                                                  
 52    |3509A               |1.2E+00               |+/-5   %     |10^-26 erg/cm^2/s/Hz|8.55E+14 |1.21E-02    |6.03E-04                  |6.03E-04                  |                           |                           |+/-6.03E-04    |Jy       |1970ApJ...162..743A|estimated error               |3509       A       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |8" aperture                             |From new raw data                                                                                                                                                  
 53    |u (SDSS) AB         |1.1E+01               |+/-0.05      |mag                 |8.44E+14 |2.10E-01    |9.70E-03                  |9.70E-03                  |                           |                           |+/-9.70E-03    |Jy       |2014ApJS..212...18B|uncertainty                   |3551   A           |Broad-band measurement                                                 |40.66969000 -0.01318000 (J2000)  |Flux in fixed aperture                                  |155"x180" aperture                      |From new raw data; Extinction-corrected for Milky Way                                                                                                              
 54    |u (SDSS) AB         |1.1E+01               |+/-0.05      |mag                 |8.44E+14 |1.71E-01    |7.88E-03                  |7.88E-03                  |                           |                           |+/-7.88E-03    |Jy       |2014ApJS..212...18B|uncertainty                   |3551   A           |Broad-band measurement                                                 |40.66969000 -0.01318000 (J2000)  |Flux in fixed aperture                                  |155"x180" aperture                      |From new raw data                                                                                                                                                  
 55    |3571A               |1.2E+00               |+/-5   %     |10^-26 erg/cm^2/s/Hz|8.40E+14 |1.22E-02    |6.12E-04                  |6.12E-04                  |                           |                           |+/-6.12E-04    |Jy       |1970ApJ...162..743A|estimated error               |3571       A       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |8" aperture                             |From new raw data                                                                                                                                                  
 56    |3636A               |1.3E+00               |+/-5   %     |10^-26 erg/cm^2/s/Hz|8.25E+14 |1.25E-02    |6.27E-04                  |6.27E-04                  |                           |                           |+/-6.27E-04    |Jy       |1970ApJ...162..743A|estimated error               |3636       A       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |8" aperture                             |From new raw data                                                                                                                                                  
 57    |U (U_T^0)           |9.5E+00               |             |mag                 |8.19E+14 |2.79E-01    |                          |                          |                           |                           |               |Jy       |1991RC3.9.C...0000d|no uncertainty reported       |3660       A       |Broad-band measurement                                                 |024006.5 -001332 (B1950)         |Multiple methods                                        |                                        |Homogenized from new and previously published data;Extinction-corrected for internal and Milky Way and K-correction applied; Standard Johnson UBVRI filters assumed
 58    |U (U_T)             |9.7E+00               |+/-0.10      |mag                 |8.19E+14 |2.39E-01    |2.31E-02                  |2.31E-02                  |                           |                           |+/-2.31E-02    |Jy       |1991RC3.9.C...0000d|rms uncertainty               |3660       A       |Broad-band measurement                                                 |024006.5 -001332 (B1950)         |Multiple methods                                        |                                        |Homogenized from new and previously published data; StandardJohnson UBVRI filters assumed                                                                          
 59    |3704A               |1.3E+00               |+/-5   %     |10^-26 erg/cm^2/s/Hz|8.10E+14 |1.27E-02    |6.34E-04                  |6.34E-04                  |                           |                           |+/-6.34E-04    |Jy       |1970ApJ...162..743A|estimated error               |3704       A       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |8" aperture                             |From new raw data                                                                                                                                                  
 62    |3862A               |1.5E+00               |+/-5   %     |10^-26 erg/cm^2/s/Hz|7.77E+14 |1.48E-02    |7.42E-04                  |7.42E-04                  |                           |                           |+/-7.42E-04    |Jy       |1970ApJ...162..743A|estimated error               |3862       A       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |8" aperture                             |From new raw data                                                                                                                                                  
 63    |4032A               |1.5E+00               |+/-5   %     |10^-26 erg/cm^2/s/Hz|7.44E+14 |1.48E-02    |7.39E-04                  |7.39E-04                  |                           |                           |+/-7.39E-04    |Jy       |1970ApJ...162..743A|estimated error               |4032       A       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |8" aperture                             |From new raw data                                                                                                                                                  
 66    |4167A               |1.5E+00               |+/-5   %     |10^-26 erg/cm^2/s/Hz|7.20E+14 |1.48E-02    |7.38E-04                  |7.38E-04                  |                           |                           |+/-7.38E-04    |Jy       |1970ApJ...162..743A|estimated error               |4167       A       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |8" aperture                             |From new raw data                                                                                                                                                  
 67    |4255A               |1.5E+00               |+/-5   %     |10^-26 erg/cm^2/s/Hz|7.05E+14 |1.54E-02    |7.72E-04                  |7.72E-04                  |                           |                           |+/-7.72E-04    |Jy       |1970ApJ...162..743A|estimated error               |4255       A       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |8" aperture                             |From new raw data                                                                                                                                                  
 68    |4250 A (OAO)        |9.0E+00               |+/-0.02      |mag                 |7.05E+14 |5.45E-01    |1.01E-02                  |1.01E-02                  |                           |                           |+/-1.01E-02    |Jy       |1982ApJ...256....1C|rms noise                     |4250       A       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |Aperture 10.0 arcmin                    |From new raw data                                                                                                                                                  
 71    |4350A               |1.7E+00               |+/-5   %     |10^-26 erg/cm^2/s/Hz|6.90E+14 |1.66E-02    |8.31E-04                  |8.31E-04                  |                           |                           |+/-8.31E-04    |Jy       |1970ApJ...162..743A|estimated error               |4350       A       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |8" aperture                             |From new raw data                                                                                                                                                  
 72    |m_p                 |9.7E+00               |+/-0.4       |mag                 |6.81E+14 |5.62E-01    |2.50E-01                  |2.50E-01                  |                           |                           |+/-2.50E-01    |Jy       |1965CGCG5.C...0000Z|rms noise                     |4400       A       |Broad-band measurement                                                 |024006.0 -001300. (B1950)        |Estimated by eye                                        |                                        |From new raw data                                                                                                                                                  
 73    |B (B_T)             |9.6E+00               |+/-0.10      |mag                 |6.81E+14 |6.10E-01    |5.89E-02                  |5.89E-02                  |                           |                           |+/-5.89E-02    |Jy       |1991RC3.9.C...0000d|rms uncertainty               |4400       A       |Broad-band measurement                                                 |024006.5 -001332 (B1950)         |Multiple methods                                        |                                        |Homogenized from new and previously published data; StandardJohnson UBVRI filters assumed                                                                          
 74    |B (m_B)             |9.7E+00               |+/-0.15      |mag                 |6.81E+14 |5.77E-01    |8.55E-02                  |8.55E-02                  |                           |                           |+/-8.55E-02    |Jy       |1991RC3.9.C...0000d|rms uncertainty               |4400       A       |Broad-band measurement                                                 |024006.5 -001332 (B1950)         |Multiple methods                                        |                                        |Homogenized from new and previously published data; StandardJohnson UBVRI filters assumed                                                                          
 75    |B (B_T^0)           |9.5E+00               |             |mag                 |6.81E+14 |6.94E-01    |                          |                          |                           |                           |               |Jy       |1991RC3.9.C...0000d|no uncertainty reported       |4400       A       |Broad-band measurement                                                 |024006.5 -001332 (B1950)         |Multiple methods                                        |                                        |Homogenized from new and previously published data;Extinction-corrected for internal and Milky Way and K-correction applied; Standard Johnson UBVRI filters assumed
 76    |4464A               |1.6E+00               |+/-5   %     |10^-26 erg/cm^2/s/Hz|6.72E+14 |1.62E-02    |8.09E-04                  |8.09E-04                  |                           |                           |+/-8.09E-04    |Jy       |1970ApJ...162..743A|estimated error               |4464       A       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |8" aperture                             |From new raw data                                                                                                                                                  
 77    |4566A               |1.7E+00               |+/-5   %     |10^-26 erg/cm^2/s/Hz|6.57E+14 |1.66E-02    |8.29E-04                  |8.29E-04                  |                           |                           |+/-8.29E-04    |Jy       |1970ApJ...162..743A|estimated error               |4566       A       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |8" aperture                             |From new raw data                                                                                                                                                  
 78    |B_J                 |1.0E+01               |             |mag                 |6.41E+14 |3.08E-01    |                          |                          |                           |                           |               |Jy       |2005MNRAS.361...34D|no uncertainty reported       |4680   A           |Broad-band measurement                                                 |024240.6 -000047.5 (J2000)       |Flux in fixed aperture                                  |                                        |From new raw data                                                                                                                                                  
 80    |g (SDSS) AB         |9.4E+00               |+/-0.05      |mag                 |6.40E+14 |6.17E-01    |2.84E-02                  |2.84E-02                  |                           |                           |+/-2.84E-02    |Jy       |2014ApJS..212...18B|uncertainty                   |4681   A           |Broad-band measurement                                                 |40.66969000 -0.01318000 (J2000)  |Flux in fixed aperture                                  |155"x180" aperture                      |From new raw data; Extinction-corrected for Milky Way                                                                                                              
 81    |g (SDSS) AB         |9.6E+00               |+/-0.05      |mag                 |6.40E+14 |5.25E-01    |2.42E-02                  |2.42E-02                  |                           |                           |+/-2.42E-02    |Jy       |2014ApJS..212...18B|uncertainty                   |4681   A           |Broad-band measurement                                                 |40.66969000 -0.01318000 (J2000)  |Flux in fixed aperture                                  |155"x180" aperture                      |From new raw data                                                                                                                                                  
 82    |4785A               |1.7E+00               |+/-5   %     |10^-26 erg/cm^2/s/Hz|6.27E+14 |1.72E-02    |8.58E-04                  |8.58E-04                  |                           |                           |+/-8.58E-04    |Jy       |1970ApJ...162..743A|estimated error               |4785       A       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |8" aperture                             |From new raw data                                                                                                                                                  
 85    |4900A               |1.8E+00               |+/-5   %     |10^-26 erg/cm^2/s/Hz|6.12E+14 |1.84E-02    |9.21E-04                  |9.21E-04                  |                           |                           |+/-9.21E-04    |Jy       |1970ApJ...162..743A|estimated error               |4900       A       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |8" aperture                             |From new raw data                                                                                                                                                  
 86    |4950A               |2.0E+00               |+/-5   %     |10^-26 erg/cm^2/s/Hz|6.06E+14 |2.05E-02    |1.02E-03                  |1.02E-03                  |                           |                           |+/-1.02E-03    |Jy       |1970ApJ...162..743A|estimated error               |4950       A       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |8" aperture                             |From new raw data                                                                                                                                                  
 87    |5000A               |2.5E+00               |+/-5   %     |10^-26 erg/cm^2/s/Hz|6.00E+14 |2.45E-02    |1.23E-03                  |1.23E-03                  |                           |                           |+/-1.23E-03    |Jy       |1970ApJ...162..743A|estimated error               |5000       A       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |8" aperture                             |From new raw data                                                                                                                                                  
 92    |5050A               |2.2E+00               |+/-5   %     |10^-26 erg/cm^2/s/Hz|5.94E+14 |2.24E-02    |1.12E-03                  |1.12E-03                  |                           |                           |+/-1.12E-03    |Jy       |1970ApJ...162..743A|estimated error               |5050       A       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |8" aperture                             |From new raw data                                                                                                                                                  
 93    |5100A               |1.8E+00               |+/-5   %     |10^-26 erg/cm^2/s/Hz|5.88E+14 |1.76E-02    |8.82E-04                  |8.82E-04                  |                           |                           |+/-8.82E-04    |Jy       |1970ApJ...162..743A|estimated error               |5100       A       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |8" aperture                             |From new raw data                                                                                                                                                  
 94    |5263A               |1.8E+00               |+/-5   %     |10^-26 erg/cm^2/s/Hz|5.70E+14 |1.80E-02    |9.00E-04                  |9.00E-04                  |                           |                           |+/-9.00E-04    |Jy       |1970ApJ...162..743A|estimated error               |5263       A       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |8" aperture                             |From new raw data                                                                                                                                                  
 95    |5350A               |1.8E+00               |+/-5   %     |10^-26 erg/cm^2/s/Hz|5.61E+14 |1.84E-02    |9.19E-04                  |9.19E-04                  |                           |                           |+/-9.19E-04    |Jy       |1970ApJ...162..743A|estimated error               |5350       A       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |8" aperture                             |From new raw data                                                                                                                                                  
 96    |V (Johnson)         |1.1E+01               |+/-0.05      |mag                 |5.42E+14 |1.42E-01    |6.71E-03                  |6.71E-03                  |                           |                           |+/-6.71E-03    |Jy       |1978ApJS...38..267O|uncertainty                   |5530   A           |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |18" aperture                            |From new raw data                                                                                                                                                  
 97    |V (Johnson)         |1.1E+01               |+/-0.05      |mag                 |5.42E+14 |1.16E-01    |5.47E-03                  |5.47E-03                  |                           |                           |+/-5.47E-03    |Jy       |1967ApJ...147..394P|uncertainty                   |5530 A             |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |15" aperture                            |From new raw data                                                                                                                                                  
 98    |V (Johnson)         |1.1E+01               |             |mag                 |5.42E+14 |1.03E-01    |                          |                          |                           |                           |               |Jy       |1973ApJ...183..711S|no uncertainty reported       |5530 A             |Broad-band measurement; photometric system transformed                 |                                 |Flux in fixed aperture                                  |7.6" aperture                           |From new raw data                                                                                                                                                  
 99    |V (Johnson)         |1.1E+01               |             |mag                 |5.42E+14 |1.52E-01    |                          |                          |                           |                           |               |Jy       |1973ApJ...183..711S|no uncertainty reported       |5530 A             |Broad-band measurement; photometric system transformed                 |                                 |Flux in fixed aperture                                  |12.2" aperture                          |From new raw data                                                                                                                                                  
 100   |V (Johnson)         |1.2E+01               |             |mag                 |5.42E+14 |7.20E-02    |                          |                          |                           |                           |               |Jy       |1973ApJ...183..711S|no uncertainty reported       |5530 A             |Broad-band measurement; photometric system transformed                 |                                 |Flux in fixed aperture                                  |4.9" aperture                           |From new raw data                                                                                                                                                  
 101   |V (Johnson)         |1.1E+01               |             |mag                 |5.42E+14 |1.71E-01    |                          |                          |                           |                           |               |Jy       |1973ApJ...183..711S|no uncertainty reported       |5530 A             |Broad-band measurement; photometric system transformed                 |                                 |Flux in fixed aperture                                  |15.2" aperture                          |From new raw data                                                                                                                                                  
 102   |V (Johnson)         |1.1E+01               |             |mag                 |5.42E+14 |1.41E-01    |                          |                          |                           |                           |               |Jy       |1973ApJ...183..711S|no uncertainty reported       |5530 A             |Broad-band measurement; photometric system transformed                 |                                 |Flux in fixed aperture                                  |11.4" aperture                          |From new raw data                                                                                                                                                  
 103   |V (V_T^0)           |8.8E+00               |             |mag                 |5.42E+14 |1.13E+00    |                          |                          |                           |                           |               |Jy       |1991RC3.9.C...0000d|no uncertainty reported       |5530       A       |Broad-band measurement                                                 |024006.5 -001332 (B1950)         |Multiple methods                                        |                                        |Homogenized from new and previously published data;Extinction-corrected for internal and Milky Way and K-correction applied; Standard Johnson UBVRI filters assumed
 104   |V (V_T)             |8.9E+00               |+/-0.10      |mag                 |5.42E+14 |1.03E+00    |1.00E-01                  |1.00E-01                  |                           |                           |+/-1.00E-01    |Jy       |1991RC3.9.C...0000d|rms uncertainty               |5530       A       |Broad-band measurement                                                 |024006.5 -001332 (B1950)         |Multiple methods                                        |                                        |Homogenized from new and previously published data; StandardJohnson UBVRI filters assumed                                                                          
 105   |5556A               |1.9E+00               |+/-5   %     |10^-26 erg/cm^2/s/Hz|5.40E+14 |1.86E-02    |9.33E-04                  |9.33E-04                  |                           |                           |+/-9.33E-04    |Jy       |1970ApJ...162..743A|estimated error               |5556       A       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |8" aperture                             |From new raw data                                                                                                                                                  
 106   |5840A               |1.9E+00               |+/-5   %     |10^-26 erg/cm^2/s/Hz|5.14E+14 |1.91E-02    |9.53E-04                  |9.53E-04                  |                           |                           |+/-9.53E-04    |Jy       |1970ApJ...162..743A|estimated error               |5840       A       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |8" aperture                             |From new raw data                                                                                                                                                  
 107   |6055A               |1.9E+00               |+/-5   %     |10^-26 erg/cm^2/s/Hz|4.95E+14 |1.93E-02    |9.67E-04                  |9.67E-04                  |                           |                           |+/-9.67E-04    |Jy       |1970ApJ...162..743A|estimated error               |6055       A       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |8" aperture                             |From new raw data                                                                                                                                                  
 109   |r (SDSS) AB         |9.0E+00               |+/-0.05      |mag                 |4.86E+14 |9.55E-01    |4.40E-02                  |4.40E-02                  |                           |                           |+/-4.40E-02    |Jy       |2014ApJS..212...18B|uncertainty                   |6165   A           |Broad-band measurement                                                 |40.66969000 -0.01318000 (J2000)  |Flux in fixed aperture                                  |155"x180" aperture                      |From new raw data                                                                                                                                                  
 110   |r (SDSS) AB         |8.8E+00               |+/-0.05      |mag                 |4.86E+14 |1.07E+00    |4.91E-02                  |4.91E-02                  |                           |                           |+/-4.91E-02    |Jy       |2014ApJS..212...18B|uncertainty                   |6165   A           |Broad-band measurement                                                 |40.66969000 -0.01318000 (J2000)  |Flux in fixed aperture                                  |155"x180" aperture                      |From new raw data; Extinction-corrected for Milky Way                                                                                                              
 113   |6370A               |2.0E+00               |+/-5   %     |10^-26 erg/cm^2/s/Hz|4.71E+14 |1.99E-02    |9.94E-04                  |9.94E-04                  |                           |                           |+/-9.94E-04    |Jy       |1970ApJ...162..743A|estimated error               |6370       A       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |8" aperture                             |From new raw data                                                                                                                                                  
 115   |R                   |1.0E+01               |             |mag                 |4.68E+14 |2.69E-01    |                          |                          |                           |                           |               |Jy       |2005MNRAS.361...34D|no uncertainty reported       |6400   A           |Broad-band measurement                                                 |024240.6 -000047.5 (J2000)       |Flux in fixed aperture                                  |                                        |From new raw data                                                                                                                                                  
 116   |6520A               |2.0E+00               |+/-5   %     |10^-26 erg/cm^2/s/Hz|4.60E+14 |1.98E-02    |9.91E-04                  |9.91E-04                  |                           |                           |+/-9.91E-04    |Jy       |1970ApJ...162..743A|estimated error               |6520       A       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |8" aperture                             |From new raw data                                                                                                                                                  
 117   |6540A               |2.1E+00               |+/-5   %     |10^-26 erg/cm^2/s/Hz|4.59E+14 |2.15E-02    |1.08E-03                  |1.08E-03                  |                           |                           |+/-1.08E-03    |Jy       |1970ApJ...162..743A|estimated error               |6540       A       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |8" aperture                             |From new raw data                                                                                                                                                  
 118   |6560A               |2.5E+00               |+/-5   %     |10^-26 erg/cm^2/s/Hz|4.57E+14 |2.49E-02    |1.25E-03                  |1.25E-03                  |                           |                           |+/-1.25E-03    |Jy       |1970ApJ...162..743A|estimated error               |6560       A       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |8" aperture                             |From new raw data                                                                                                                                                  
 120   |6580A               |2.7E+00               |+/-5   %     |10^-26 erg/cm^2/s/Hz|4.56E+14 |2.71E-02    |1.36E-03                  |1.36E-03                  |                           |                           |+/-1.36E-03    |Jy       |1970ApJ...162..743A|estimated error               |6580       A       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |8" aperture                             |From new raw data                                                                                                                                                  
 121   |6600A               |2.7E+00               |+/-5   %     |10^-26 erg/cm^2/s/Hz|4.55E+14 |2.75E-02    |1.37E-03                  |1.37E-03                  |                           |                           |+/-1.37E-03    |Jy       |1970ApJ...162..743A|estimated error               |6600       A       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |8" aperture                             |From new raw data                                                                                                                                                  
 123   |6620A               |2.6E+00               |+/-5   %     |10^-26 erg/cm^2/s/Hz|4.53E+14 |2.59E-02    |1.30E-03                  |1.30E-03                  |                           |                           |+/-1.30E-03    |Jy       |1970ApJ...162..743A|estimated error               |6620       A       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |8" aperture                             |From new raw data                                                                                                                                                  
 124   |6640A               |2.2E+00               |+/-5   %     |10^-26 erg/cm^2/s/Hz|4.52E+14 |2.15E-02    |1.08E-03                  |1.08E-03                  |                           |                           |+/-1.08E-03    |Jy       |1970ApJ...162..743A|estimated error               |6640       A       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |8" aperture                             |From new raw data                                                                                                                                                  
 125   |6726A               |2.2E+00               |+/-5   %     |10^-26 erg/cm^2/s/Hz|4.46E+14 |2.16E-02    |1.08E-03                  |1.08E-03                  |                           |                           |+/-1.08E-03    |Jy       |1970ApJ...162..743A|estimated error               |6726       A       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |8" aperture                             |From new raw data                                                                                                                                                  
 128   |6800A               |2.0E+00               |+/-5   %     |10^-26 erg/cm^2/s/Hz|4.41E+14 |2.00E-02    |1.00E-03                  |1.00E-03                  |                           |                           |+/-1.00E-03    |Jy       |1970ApJ...162..743A|estimated error               |6800       A       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |8" aperture                             |From new raw data                                                                                                                                                  
 129   |R (Johnson)         |1.0E+01               |+/-0.05      |mag                 |4.28E+14 |1.77E-01    |8.34E-03                  |8.34E-03                  |                           |                           |+/-8.34E-03    |Jy       |1967ApJ...147..394P|uncertainty                   |7000 A             |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |15" aperture                            |From new raw data                                                                                                                                                  
 130   |R (Johnson)         |1.0E+01               |             |mag                 |4.28E+14 |2.73E-01    |                          |                          |                           |                           |               |Jy       |1973ApJ...183..711S|no uncertainty reported       |7000 A             |Broad-band measurement; photometric system transformed                 |                                 |Flux in fixed aperture                                  |15.2" aperture                          |From new raw data; derived from a flux in a different bandand a color                                                                                              
 131   |R (Johnson)         |1.0E+01               |             |mag                 |4.28E+14 |2.27E-01    |                          |                          |                           |                           |               |Jy       |1973ApJ...183..711S|no uncertainty reported       |7000 A             |Broad-band measurement; photometric system transformed                 |                                 |Flux in fixed aperture                                  |12.2" aperture                          |From new raw data; derived from a flux in a different bandand a color                                                                                              
 132   |R (Johnson)         |1.1E+01               |             |mag                 |4.28E+14 |1.49E-01    |                          |                          |                           |                           |               |Jy       |1973ApJ...183..711S|no uncertainty reported       |7000 A             |Broad-band measurement; photometric system transformed                 |                                 |Flux in fixed aperture                                  |7.6" aperture                           |From new raw data; derived from a flux in a different bandand a color                                                                                              
 133   |R (Johnson)         |1.0E+01               |+/-0.05      |mag                 |4.28E+14 |2.17E-01    |1.02E-02                  |1.02E-02                  |                           |                           |+/-1.02E-02    |Jy       |1978ApJS...38..267O|uncertainty                   |7000   A           |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |18" aperture                            |From new raw data                                                                                                                                                  
 134   |R (Johnson)         |1.1E+01               |             |mag                 |4.28E+14 |9.55E-02    |                          |                          |                           |                           |               |Jy       |1973ApJ...183..711S|no uncertainty reported       |7000 A             |Broad-band measurement; photometric system transformed                 |                                 |Flux in fixed aperture                                  |4.9" aperture                           |From new raw data; derived from a flux in a different bandand a color                                                                                              
 135   |R (Johnson)         |1.0E+01               |             |mag                 |4.28E+14 |2.21E-01    |                          |                          |                           |                           |               |Jy       |1973ApJ...183..711S|no uncertainty reported       |7000 A             |Broad-band measurement; photometric system transformed                 |                                 |Flux in fixed aperture                                  |11.4" aperture                          |From new raw data; derived from a flux in a different bandand a color                                                                                              
 136   |7100A               |2.0E+00               |+/-5   %     |10^-26 erg/cm^2/s/Hz|4.23E+14 |2.04E-02    |1.02E-03                  |1.02E-03                  |                           |                           |+/-1.02E-03    |Jy       |1970ApJ...162..743A|estimated error               |7100       A       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |8" aperture                             |From new raw data                                                                                                                                                  
 137   |i (SDSS) AB         |8.5E+00               |+/-0.05      |mag                 |4.01E+14 |1.41E+00    |6.48E-02                  |6.48E-02                  |                           |                           |+/-6.48E-02    |Jy       |2014ApJS..212...18B|uncertainty                   |7480   A           |Broad-band measurement                                                 |40.66969000 -0.01318000 (J2000)  |Flux in fixed aperture                                  |155"x180" aperture                      |From new raw data; Extinction-corrected for Milky Way                                                                                                              
 138   |i (SDSS) AB         |8.6E+00               |+/-0.05      |mag                 |4.01E+14 |1.30E+00    |5.96E-02                  |5.96E-02                  |                           |                           |+/-5.96E-02    |Jy       |2014ApJS..212...18B|uncertainty                   |7480   A           |Broad-band measurement                                                 |40.66969000 -0.01318000 (J2000)  |Flux in fixed aperture                                  |155"x180" aperture                      |From new raw data                                                                                                                                                  
 139   |7530A               |2.1E+00               |+/-5   %     |10^-26 erg/cm^2/s/Hz|3.98E+14 |2.09E-02    |1.04E-03                  |1.04E-03                  |                           |                           |+/-1.04E-03    |Jy       |1970ApJ...162..743A|estimated error               |7530       A       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |8" aperture                             |From new raw data                                                                                                                                                  
 140   |7850A               |2.1E+00               |+/-5   %     |10^-26 erg/cm^2/s/Hz|3.82E+14 |2.12E-02    |1.06E-03                  |1.06E-03                  |                           |                           |+/-1.06E-03    |Jy       |1970ApJ...162..743A|estimated error               |7850       A       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |8" aperture                             |From new raw data                                                                                                                                                  
 142   |I                   |9.9E+00               |             |mag                 |3.79E+14 |2.79E-01    |                          |                          |                           |                           |               |Jy       |2005MNRAS.361...34D|no uncertainty reported       |7900   A           |Broad-band measurement                                                 |024240.6 -000047.5 (J2000)       |Flux in fixed aperture                                  |                                        |From new raw data                                                                                                                                                  
 143   |8080A               |2.1E+00               |+/-10  %     |10^-26 erg/cm^2/s/Hz|3.71E+14 |2.13E-02    |2.13E-03                  |2.13E-03                  |                           |                           |+/-2.13E-03    |Jy       |1970ApJ...162..743A|estimated error               |8080       A       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |8" aperture                             |From new raw data                                                                                                                                                  
 144   |8400A               |2.2E+00               |+/-10  %     |10^-26 erg/cm^2/s/Hz|3.57E+14 |2.17E-02    |2.17E-03                  |2.17E-03                  |                           |                           |+/-2.17E-03    |Jy       |1970ApJ...162..743A|estimated error               |8400       A       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |8" aperture                             |From new raw data                                                                                                                                                  
 145   |z (SDSS) AB         |8.4E+00               |+/-0.05      |mag                 |3.36E+14 |1.65E+00    |7.60E-02                  |7.60E-02                  |                           |                           |+/-7.60E-02    |Jy       |2014ApJS..212...18B|uncertainty                   |8931   A           |Broad-band measurement                                                 |40.66969000 -0.01318000 (J2000)  |Flux in fixed aperture                                  |155"x180" aperture                      |From new raw data                                                                                                                                                  
 146   |z (SDSS) AB         |8.3E+00               |+/-0.05      |mag                 |3.36E+14 |1.76E+00    |8.09E-02                  |8.09E-02                  |                           |                           |+/-8.09E-02    |Jy       |2014ApJS..212...18B|uncertainty                   |8931   A           |Broad-band measurement                                                 |40.66969000 -0.01318000 (J2000)  |Flux in fixed aperture                                  |155"x180" aperture                      |From new raw data; Extinction-corrected for Milky Way                                                                                                              
 147   |I (Johnson)         |9.9E+00               |+/-0.05      |mag                 |3.33E+14 |2.55E-01    |1.20E-02                  |1.20E-02                  |                           |                           |+/-1.20E-02    |Jy       |1967ApJ...147..394P|uncertainty                   |9000 A             |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |15" aperture                            |From new raw data                                                                                                                                                  
 157   |J (ESO/SPM)         |5.6E+02               |+/-37.35     |milliJy             |2.50E+14 |5.61E-01    |3.73E-02                  |3.73E-02                  |                           |                           |+/-3.73E-02    |Jy       |1995ApJ...453..616S|rms uncertainty               |1.198      microns |Broad-band measurement                                                 |024007.7 -001329 (B1950)         |Flux in fixed aperture                                  |15" aperture                            |From new raw data                                                                                                                                                  
 158   |J (RGO)             |9.1E+00               |+/-0.03      |mag                 |2.50E+14 |3.72E-01    |1.04E-02                  |1.04E-02                  |                           |                           |+/-1.04E-02    |Jy       |1981MNRAS.197.1067G|uncertainty                   |1.20    microns    |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |12" aperture                            |From new raw data                                                                                                                                                  
 159   |J (2MASS) AB        |7.9E+00               |+/-0.05      |mag                 |2.43E+14 |2.63E+00    |1.21E-01                  |1.21E-01                  |                           |                           |+/-1.21E-01    |Jy       |2014ApJS..212...18B|uncertainty                   |12320   A          |Broad-band measurement                                                 |40.66969000 -0.01318000 (J2000)  |Flux in fixed aperture                                  |155"x180" aperture                      |From new raw data; Extinction-corrected for Milky Way                                                                                                              
 160   |J (2MASS) AB        |7.9E+00               |+/-0.05      |mag                 |2.43E+14 |2.54E+00    |1.17E-01                  |1.17E-01                  |                           |                           |+/-1.17E-01    |Jy       |2014ApJS..212...18B|uncertainty                   |12320   A          |Broad-band measurement                                                 |40.66969000 -0.01318000 (J2000)  |Flux in fixed aperture                                  |155"x180" aperture                      |From new raw data                                                                                                                                                  
 161   |J (Johnson)         |7.6E+00               |+/-0.03      |mag                 |2.42E+14 |1.44E+00    |4.02E-02                  |4.02E-02                  |                           |                           |+/-4.02E-02    |Jy       |1977HarvU.T00M....A|uncertainty                   |1.24    microns    |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |53.4" aperture                          |From new raw data; derived from a flux in a different bandand a color                                                                                              
 162   |J (Johnson)         |7.2E+00               |+/-0.03      |mag                 |2.42E+14 |2.09E+00    |5.87E-02                  |5.87E-02                  |                           |                           |+/-5.87E-02    |Jy       |1977HarvU.T00M....A|uncertainty                   |1.24    microns    |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |105" aperture                           |From new raw data; derived from a flux in a different bandand a color                                                                                              
 163   |J (Johnson)         |8.1E+00               |+/-0.03      |mag                 |2.42E+14 |8.89E-01    |2.49E-02                  |2.49E-02                  |                           |                           |+/-2.49E-02    |Jy       |1977HarvU.T00M....A|uncertainty                   |1.24    microns    |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |27.4" aperture                          |From new raw data; derived from a flux in a different bandand a color                                                                                              
 164   |F_J (total)         |3.6E+00               |+/-3.02      |log milliJy         |2.41E+14 |4.07E+00    |1.05E+00                  |1.05E+00                  |                           |                           |+/-1.05E+00    |Jy       |1995ApJ...453..616S|1 sigma                       |1.244      microns |Broad-band measurement                                                 |                                 |Corrected to total flux from single aperture measurement|                                        |Homogenized from new and previously published data                                                                                                                 
 165   |J_20 (2MASS LGA)    |7.0E+00               |+/-0.015     |mag                 |2.40E+14 |2.49E+00    |3.47E-02                  |3.47E-02                  |                           |                           |+/-3.47E-02    |Jy       |2003AJ....125..525J|1 sigma uncert.               |1.25      microns  |Broad-band measurement                                                 |024240.77 -000047.5 (J2000)      |Flux integrated from map                                |190.0 x  155.8 arcsec integration area. |From new raw data; Corrected for contaminating sources                                                                                                             
 166   |J_Kron (2MASS LGA)  |7.1E+00               |+/-0.015     |mag                 |2.40E+14 |2.25E+00    |3.13E-02                  |3.13E-02                  |                           |                           |+/-3.13E-02    |Jy       |2003AJ....125..525J|1 sigma uncert.               |1.25      microns  |Broad-band measurement                                                 |024240.77 -000047.5 (J2000)      |Flux integrated from map                                |127.4 x  104.5 arcsec integration area. |From new raw data; Corrected for contaminating sources                                                                                                             
 167   |J_tot (2MASS LGA)   |7.0E+00               |+/-0.015     |mag                 |2.40E+14 |2.60E+00    |3.62E-02                  |3.62E-02                  |                           |                           |+/-3.62E-02    |Jy       |2003AJ....125..525J|1 sigma uncert.               |1.25      microns  |Broad-band measurement                                                 |024240.77 -000047.5 (J2000)      |Total flux                                              |                                        |From new raw data                                                                                                                                                  
 168   |J_14arcsec (2MASS)  |8.7E+00               |+/-0.015     |mag                 |2.40E+14 |5.11E-01    |7.11E-03                  |7.11E-03                  |                           |                           |+/-7.11E-03    |Jy       |20032MASX.C.......:|1 sigma uncert.               |1.25      microns  |Broad-band measurement                                                 |024240.77 -000047.5 (J2000)      |Flux in fixed aperture                                  |14.0 x 14.0 arcsec aperture             |From new raw data                                                                                                                                                  
 169   |1.25 microns        |2.6E-01               |+/-10  %     |Jy                  |2.40E+14 |2.60E-01    |2.61E-02                  |2.61E-02                  |                           |                           |+/-2.61E-02    |Jy       |1978ApJ...226..550R|uncertainty                   |1.25    microns    |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |8.5" aperture                           |From new raw data                                                                                                                                                  
 172   |J (Johnson)         |8.8E+00               |+/-0.1       |mag                 |2.38E+14 |4.98E-01    |4.80E-02                  |4.80E-02                  |                           |                           |+/-4.80E-02    |Jy       |1967ApJ...147..394P|uncertainty                   |1.26 microns       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |15" aperture                            |From new raw data                                                                                                                                                  
 174   |J (VLT)             |                      |<0.0084      |Jy                  |2.30E+14 |            |                          |                          |0.00840000                 |                           |<8.40E-03      |Jy       |2008A&A...485...33H|no uncertainty reported       |1.3 microns        |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |Nuclear flux                            |From new raw data                                                                                                                                                  
 176   |H' (Johnson)        |8.2E+00               |             |mag                 |1.93E+14 |6.71E-01    |                          |                          |                           |                           |               |Jy       |1968AJ.....73..866W|no uncertainty reported       |1.55 microns       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |13" aperture;Low quality data           |Averaged from previously published data                                                                                                                            
 177   |H' (Johnson)        |9.1E+00               |             |mag                 |1.93E+14 |2.82E-01    |                          |                          |                           |                           |               |Jy       |1968AJ.....73..866W|no uncertainty reported       |1.55 microns       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |13" aperture;Low quality data           |Averaged from previously published data                                                                                                                            
 178   |H (ESO/SPM)         |7.7E+02               |+/-51.49     |milliJy             |1.90E+14 |7.73E-01    |5.15E-02                  |5.15E-02                  |                           |                           |+/-5.15E-02    |Jy       |1995ApJ...453..616S|rms uncertainty               |1.580      microns |Broad-band measurement                                                 |024007.7 -001329 (B1950)         |Flux in fixed aperture                                  |15" aperture                            |From new raw data                                                                                                                                                  
 179   |H (Johnson)         |7.9E+00               |+/-0.1       |mag                 |1.85E+14 |8.18E-01    |7.89E-02                  |7.89E-02                  |                           |                           |+/-7.89E-02    |Jy       |1967ApJ...147..394P|uncertainty                   |1.62 microns       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |15" aperture                            |From new raw data                                                                                                                                                  
 180   |F_H (total)         |3.8E+00               |+/-3.18      |log milliJy         |1.84E+14 |5.89E+00    |1.52E+00                  |1.52E+00                  |                           |                           |+/-1.52E+00    |Jy       |1995ApJ...453..616S|1 sigma                       |1.634      microns |Broad-band measurement                                                 |                                 |Corrected to total flux from single aperture measurement|                                        |Homogenized from new and previously published data                                                                                                                 
 181   |1.6 microns         |3.5E-01               |+/-10  %     |Jy                  |1.84E+14 |3.50E-01    |3.54E-02                  |3.54E-02                  |                           |                           |+/-3.54E-02    |Jy       |1978ApJ...226..550R|uncertainty                   |1.63    microns    |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |8.5" aperture                           |From new raw data                                                                                                                                                  
 182   |H (RGO)             |8.2E+00               |+/-0.03      |mag                 |1.83E+14 |5.31E-01    |1.49E-02                  |1.49E-02                  |                           |                           |+/-1.49E-02    |Jy       |1981MNRAS.197.1067G|uncertainty                   |1.64    microns    |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |12" aperture                            |From new raw data                                                                                                                                                  
 183   |H_20 (2MASS LGA)    |6.3E+00               |+/-0.015     |mag                 |1.82E+14 |3.13E+00    |4.36E-02                  |4.36E-02                  |                           |                           |+/-4.36E-02    |Jy       |2003AJ....125..525J|1 sigma uncert.               |1.65      microns  |Broad-band measurement                                                 |024240.77 -000047.5 (J2000)      |Flux integrated from map                                |190.0 x  155.8 arcsec integration area. |From new raw data; Corrected for contaminating sources                                                                                                             
 184   |H_Kron (2MASS LGA)  |6.4E+00               |+/-0.015     |mag                 |1.82E+14 |2.88E+00    |4.01E-02                  |4.01E-02                  |                           |                           |+/-4.01E-02    |Jy       |2003AJ....125..525J|1 sigma uncert.               |1.65      microns  |Broad-band measurement                                                 |024240.77 -000047.5 (J2000)      |Flux integrated from map                                |127.4 x  104.5 arcsec integration area. |From new raw data; Corrected for contaminating sources                                                                                                             
 185   |H_tot (2MASS LGA)   |6.3E+00               |+/-0.015     |mag                 |1.82E+14 |3.21E+00    |4.47E-02                  |4.47E-02                  |                           |                           |+/-4.47E-02    |Jy       |2003AJ....125..525J|1 sigma uncert.               |1.65      microns  |Broad-band measurement                                                 |024240.77 -000047.5 (J2000)      |Total flux                                              |                                        |From new raw data                                                                                                                                                  
 186   |H_14arcsec (2MASS)  |7.9E+00               |+/-0.015     |mag                 |1.82E+14 |7.34E-01    |1.02E-02                  |1.02E-02                  |                           |                           |+/-1.02E-02    |Jy       |20032MASX.C.......:|1 sigma uncert.               |1.65      microns  |Broad-band measurement                                                 |024240.77 -000047.5 (J2000)      |Flux in fixed aperture                                  |14.0 x 14.0 arcsec aperture             |From new raw data                                                                                                                                                  
 188   |H (2MASS) AB        |7.6E+00               |+/-0.05      |mag                 |1.82E+14 |3.24E+00    |1.49E-01                  |1.49E-01                  |                           |                           |+/-1.49E-01    |Jy       |2014ApJS..212...18B|uncertainty                   |16440   A          |Broad-band measurement                                                 |40.66969000 -0.01318000 (J2000)  |Flux in fixed aperture                                  |155"x180" aperture                      |From new raw data; Extinction-corrected for Milky Way                                                                                                              
 189   |H (2MASS) AB        |7.7E+00               |+/-0.05      |mag                 |1.82E+14 |3.17E+00    |1.46E-01                  |1.46E-01                  |                           |                           |+/-1.46E-01    |Jy       |2014ApJS..212...18B|uncertainty                   |16440   A          |Broad-band measurement                                                 |40.66969000 -0.01318000 (J2000)  |Flux in fixed aperture                                  |155"x180" aperture                      |From new raw data                                                                                                                                                  
 190   |H                   |7.9E+00               |+/-0.06      |mag                 |1.82E+14 |6.85E-01    |3.89E-02                  |3.89E-02                  |                           |                           |+/-3.89E-02    |Jy       |1978ApJS...38..267O|uncertainty                   |1.65    microns    |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |18" aperture                            |Averaged new and previously published data                                                                                                                         
 191   |H                   |8.5E+00               |+/-0.06      |mag                 |1.82E+14 |4.02E-01    |2.28E-02                  |2.28E-02                  |                           |                           |+/-2.28E-02    |Jy       |1978ApJS...38..267O|uncertainty                   |1.65    microns    |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |9" aperture                             |Averaged new and previously published data                                                                                                                         
 192   |1.6 microns         |8.0E+00               |             |mag                 |1.82E+14 |6.30E-01    |                          |                          |                           |                           |               |Jy       |1974MNRAS.169..357P|no uncertainty reported       |1.65   microns     |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |13.5" aperture                          |Averaged new and previously published data                                                                                                                         
 193   |1.6 microns         |7.4E+00               |             |mag                 |1.82E+14 |1.12E+00    |                          |                          |                           |                           |               |Jy       |1974MNRAS.169..357P|no uncertainty reported       |1.65   microns     |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |32" aperture                            |Averaged new and previously published data                                                                                                                         
 194   |1.6 microns         |8.5E+00               |+/-0.07      |mag                 |1.82E+14 |3.94E-01    |2.62E-02                  |2.62E-02                  |                           |                           |+/-2.62E-02    |Jy       |1974MNRAS.169..357P|uncertainty                   |1.65   microns     |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |10.0" aperture;Low quality data         |From new raw data                                                                                                                                                  
 195   |1.6 microns         |7.5E+00               |+/-0.10      |mag                 |1.82E+14 |9.45E-01    |9.11E-02                  |9.11E-02                  |                           |                           |+/-9.11E-02    |Jy       |1974MNRAS.169..357P|uncertainty                   |1.65   microns     |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |25" aperture                            |From new raw data                                                                                                                                                  
 196   |1.6 microns         |7.6E+00               |+/-0.10      |mag                 |1.82E+14 |9.36E-01    |9.03E-02                  |9.03E-02                  |                           |                           |+/-9.03E-02    |Jy       |1974MNRAS.169..357P|uncertainty                   |1.65   microns     |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |22" aperture;Low quality data           |From new raw data                                                                                                                                                  
 197   |1.6 microns         |7.4E+00               |             |mag                 |1.82E+14 |1.12E+00    |                          |                          |                           |                           |               |Jy       |1974MNRAS.169..357P|no uncertainty reported       |1.65   microns     |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |28" aperture                            |Averaged new and previously published data                                                                                                                         
 198   |H (Johnson)         |7.3E+00               |+/-0.03      |mag                 |1.82E+14 |1.26E+00    |3.52E-02                  |3.52E-02                  |                           |                           |+/-3.52E-02    |Jy       |1977HarvU.T00M....A|uncertainty                   |1.65    microns    |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |27.4" aperture                          |From new raw data; derived from a flux in a different bandand a color                                                                                              
 199   |1.6 microns         |7.9E+00               |             |mag                 |1.82E+14 |7.10E-01    |                          |                          |                           |                           |               |Jy       |1974MNRAS.169..357P|no uncertainty reported       |1.65   microns     |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |15" aperture                            |Averaged new and previously published data                                                                                                                         
 200   |H (Johnson)         |6.8E+00               |+/-0.03      |mag                 |1.82E+14 |2.05E+00    |5.74E-02                  |5.74E-02                  |                           |                           |+/-5.74E-02    |Jy       |1977HarvU.T00M....A|uncertainty                   |1.65    microns    |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |53.4" aperture                          |From new raw data; derived from a flux in a different bandand a color                                                                                              
 201   |H (Johnson)         |6.5E+00               |+/-0.03      |mag                 |1.82E+14 |2.83E+00    |7.92E-02                  |7.92E-02                  |                           |                           |+/-7.92E-02    |Jy       |1977HarvU.T00M....A|uncertainty                   |1.65    microns    |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |105" aperture                           |From new raw data; derived from a flux in a different bandand a color                                                                                              
 202   |H (VLT)             |2.2E-02               |             |Jy                  |1.80E+14 |2.20E-02    |                          |                          |                           |                           |               |Jy       |2008A&A...485...33H|no uncertainty reported       |1.65 microns       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |Nuclear flux                            |From new raw data                                                                                                                                                  
 208   |K (VLT)             |9.8E-02               |             |Jy                  |1.40E+14 |9.80E-02    |                          |                          |                           |                           |               |Jy       |2008A&A...485...33H|no uncertainty reported       |2.2  microns       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |Nuclear flux                            |From new raw data                                                                                                                                                  
 210   |Ks (2MASS) AB       |7.6E+00               |+/-0.05      |mag                 |1.39E+14 |3.24E+00    |1.49E-01                  |1.49E-01                  |                           |                           |+/-1.49E-01    |Jy       |2014ApJS..212...18B|uncertainty                   |21590   A          |Broad-band measurement                                                 |40.66969000 -0.01318000 (J2000)  |Flux in fixed aperture                                  |155"x180" aperture                      |From new raw data; Extinction-corrected for Milky Way                                                                                                              
 211   |Ks (2MASS) AB       |7.6E+00               |+/-0.05      |mag                 |1.39E+14 |3.19E+00    |1.47E-01                  |1.47E-01                  |                           |                           |+/-1.47E-01    |Jy       |2014ApJS..212...18B|uncertainty                   |21590   A          |Broad-band measurement                                                 |40.66969000 -0.01318000 (J2000)  |Flux in fixed aperture                                  |155"x180" aperture                      |From new raw data                                                                                                                                                  
 212   |K_20 (2MASS LGA)    |5.8E+00               |+/-0.015     |mag                 |1.38E+14 |3.16E+00    |4.39E-02                  |4.39E-02                  |                           |                           |+/-4.39E-02    |Jy       |2003AJ....125..525J|1 sigma uncert.               |2.17      microns  |Broad-band measurement                                                 |024240.77 -000047.5 (J2000)      |Flux integrated from map                                |190.0 x  155.8 arcsec integration area. |From new raw data; Corrected for contaminating sources                                                                                                             
 213   |K_Kron (2MASS LGA)  |5.9E+00               |+/-0.015     |mag                 |1.38E+14 |2.95E+00    |4.11E-02                  |4.11E-02                  |                           |                           |+/-4.11E-02    |Jy       |2003AJ....125..525J|1 sigma uncert.               |2.17      microns  |Broad-band measurement                                                 |024240.77 -000047.5 (J2000)      |Flux integrated from map                                |127.4 x  104.5 arcsec integration area. |From new raw data; Corrected for contaminating sources                                                                                                             
 214   |K_tot (2MASS LGA)   |5.8E+00               |+/-0.016     |mag                 |1.38E+14 |3.23E+00    |4.79E-02                  |4.79E-02                  |                           |                           |+/-4.79E-02    |Jy       |2003AJ....125..525J|1 sigma uncert.               |2.17      microns  |Broad-band measurement                                                 |024240.77 -000047.5 (J2000)      |Total flux                                              |                                        |From new raw data                                                                                                                                                  
 215   |K_s_14arcsec (2MASS)|7.0E+00               |+/-0.015     |mag                 |1.38E+14 |1.06E+00    |1.48E-02                  |1.48E-02                  |                           |                           |+/-1.48E-02    |Jy       |20032MASX.C.......:|1 sigma uncert.               |2.17      microns  |Broad-band measurement                                                 |024240.77 -000047.5 (J2000)      |Flux in fixed aperture                                  |14.0 x 14.0 arcsec aperture             |From new raw data                                                                                                                                                  
 216   |K_s (VLT/NACO)      |8.9E+00               |             |mag                 |1.38E+14 |1.84E-01    |                          |                          |                           |                           |               |Jy       |2006A&A...446..813G|no uncertainty reported       |2.18   microns     |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |Nuclear; aperture radius = 0.27"        |From reprocessed raw data                                                                                                                                          
 217   |K_s (VLT/NACO)      |9.3E+00               |             |mag                 |1.38E+14 |1.27E-01    |                          |                          |                           |                           |               |Jy       |2006A&A...446..813G|no uncertainty reported       |2.18   microns     |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |Nuclear; aperture radius = 0.13"        |From reprocessed raw data                                                                                                                                          
 218   |K_s (VLT/NACO)      |9.9E+00               |             |mag                 |1.38E+14 |7.31E-02    |                          |                          |                           |                           |               |Jy       |2006A&A...446..813G|no uncertainty reported       |2.18   microns     |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |Nuclear; aperture radius = 0.08"        |From reprocessed raw data                                                                                                                                          
 219   |K_s (2MASS)         |6.8E+00               |             |mag                 |1.38E+14 |1.27E+00    |                          |                          |                           |                           |               |Jy       |2006A&A...453..863P|no uncertainty reported       |2.17   microns     |Broad-band measurement                                                 |                                 |Modelled datum                                          |Disk magnitude                          |From reprocessed raw data                                                                                                                                          
 220   |K_s (2MASS)         |8.0E+00               |             |mag                 |1.38E+14 |4.13E-01    |                          |                          |                           |                           |               |Jy       |2006A&A...453..863P|no uncertainty reported       |2.17   microns     |Broad-band measurement                                                 |                                 |Modelled datum                                          |AGN magnitude                           |From reprocessed raw data                                                                                                                                          
 221   |K_s (2MASS)         |7.3E+00               |             |mag                 |1.38E+14 |7.87E-01    |                          |                          |                           |                           |               |Jy       |2006A&A...453..863P|no uncertainty reported       |2.17   microns     |Broad-band measurement                                                 |                                 |Modelled datum                                          |Bulge magnitude                         |From reprocessed raw data                                                                                                                                          
 222   |K (VLTI)            |1.3E+02               |+/-60        |milliJy             |1.38E+14 |1.30E-01    |6.00E-02                  |6.00E-02                  |                           |                           |+/-6.00E-02    |Jy       |2004A&A...418L..39W|uncertainty                   |2.18   microns     |Broad-band measurement                                                 |                                 |From fitting to map                                     |Nuclear flux; lower limit               |From new raw data                                                                                                                                                  
 224   |F_K (total)         |3.8E+00               |+/-3.25      |log milliJy         |1.37E+14 |6.92E+00    |1.79E+00                  |1.79E+00                  |                           |                           |+/-1.79E+00    |Jy       |1995ApJ...453..616S|1 sigma                       |2.194      microns |Broad-band measurement                                                 |                                 |Corrected to total flux from single aperture measurement|                                        |Homogenized from new and previously published data                                                                                                                 
 225   |K (RGO)             |7.5E+00               |+/-0.03      |mag                 |1.37E+14 |6.68E-01    |1.87E-02                  |1.87E-02                  |                           |                           |+/-1.87E-02    |Jy       |1981MNRAS.197.1067G|uncertainty                   |2.19    microns    |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |12" aperture                            |From new raw data                                                                                                                                                  
 226   |2.2 microns         |7.6E+00               |             |mag                 |1.36E+14 |5.76E-01    |                          |                          |                           |                           |               |Jy       |1974MNRAS.169..357P|no uncertainty reported       |2.2   microns      |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |10.0" aperture                          |Averaged new and previously published data                                                                                                                         
 227   |2.2 microns         |3.7E-01               |+/-0.02      |Jy                  |1.36E+14 |3.70E-01    |2.00E-02                  |2.00E-02                  |                           |                           |+/-2.00E-02    |Jy       |1972ApJ...176L..95R|1 sigma                       |2.2 microns        |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |6" aperture                             |From new raw data                                                                                                                                                  
 228   |2.2 microns         |6.8E+00               |             |mag                 |1.36E+14 |1.16E+00    |                          |                          |                           |                           |               |Jy       |1974MNRAS.169..357P|no uncertainty reported       |2.2   microns      |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |28" aperture                            |Averaged new and previously published data                                                                                                                         
 229   |2.2 microns         |6.8E+00               |             |mag                 |1.36E+14 |1.17E+00    |                          |                          |                           |                           |               |Jy       |1974MNRAS.169..357P|no uncertainty reported       |2.2   microns      |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |32" aperture                            |Averaged new and previously published data                                                                                                                         
 230   |2.2 microns         |7.3E+00               |             |mag                 |1.36E+14 |7.32E-01    |                          |                          |                           |                           |               |Jy       |1974MNRAS.169..357P|no uncertainty reported       |2.2   microns      |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |13.5" aperture                          |Averaged new and previously published data                                                                                                                         
 231   |2.2 microns         |7.1E+00               |+/-0.10      |mag                 |1.36E+14 |9.38E-01    |9.05E-02                  |9.05E-02                  |                           |                           |+/-9.05E-02    |Jy       |1974MNRAS.169..357P|uncertainty                   |2.2   microns      |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |22" aperture;Low quality data           |From new raw data                                                                                                                                                  
 232   |2.2 microns         |7.1E+00               |             |mag                 |1.36E+14 |9.13E-01    |                          |                          |                           |                           |               |Jy       |1974MNRAS.169..357P|no uncertainty reported       |2.2   microns      |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |20" aperture                            |Averaged new and previously published data                                                                                                                         
 233   |2.2 microns         |7.3E+00               |             |mag                 |1.36E+14 |7.81E-01    |                          |                          |                           |                           |               |Jy       |1974MNRAS.169..357P|no uncertainty reported       |2.2   microns      |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |15" aperture                            |Averaged new and previously published data                                                                                                                         
 234   |2.2 microns         |6.9E+00               |+/-0.10      |mag                 |1.36E+14 |1.04E+00    |1.00E-01                  |1.00E-01                  |                           |                           |+/-1.00E-01    |Jy       |1974MNRAS.169..357P|uncertainty                   |2.2   microns      |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |25" aperture;Low quality data           |From new raw data                                                                                                                                                  
 235   |K (ESO/SPM)         |9.3E+02               |+/-62.11     |milliJy             |1.36E+14 |9.33E-01    |6.21E-02                  |6.21E-02                  |                           |                           |+/-6.21E-02    |Jy       |1995ApJ...453..616S|rms uncertainty               |2.210      microns |Broad-band measurement                                                 |024007.7 -001329 (B1950)         |Flux in fixed aperture                                  |15" aperture                            |From new raw data                                                                                                                                                  
 236   |K (Johnson)         |7.2E+00               |+/-0.1       |mag                 |1.35E+14 |8.63E-01    |8.33E-02                  |8.33E-02                  |                           |                           |+/-8.33E-02    |Jy       |1967ApJ...147..394P|uncertainty                   |2.22 microns       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |15" aperture                            |From new raw data                                                                                                                                                  
 237   |2.2 microns         |5.4E-01               |+/-10  %     |Jy                  |1.35E+14 |5.40E-01    |5.40E-02                  |5.40E-02                  |                           |                           |+/-5.40E-02    |Jy       |1978ApJ...226..550R|uncertainty                   |2.22    microns    |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |8.5" aperture                           |From new raw data                                                                                                                                                  
 238   |K (Johnson)         |6.8E+00               |+/-0.03      |mag                 |1.35E+14 |1.27E+00    |3.56E-02                  |3.56E-02                  |                           |                           |+/-3.56E-02    |Jy       |1977HarvU.T00M....A|uncertainty                   |2.22    microns    |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |27.4" aperture                          |From new raw data                                                                                                                                                  
 239   |K (Johnson)         |6.1E+00               |+/-0.03      |mag                 |1.35E+14 |2.54E+00    |7.11E-02                  |7.11E-02                  |                           |                           |+/-7.11E-02    |Jy       |1977HarvU.T00M....A|uncertainty                   |2.22    microns    |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |105" aperture                           |From new raw data                                                                                                                                                  
 240   |K (Johnson)         |6.3E+00               |+/-0.03      |mag                 |1.35E+14 |1.94E+00    |5.44E-02                  |5.44E-02                  |                           |                           |+/-5.44E-02    |Jy       |1977HarvU.T00M....A|uncertainty                   |2.22    microns    |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |53.4" aperture                          |From new raw data                                                                                                                                                  
 241   |K                   |7.6E+00               |+/-0.04      |mag                 |1.31E+14 |5.43E-01    |2.04E-02                  |2.04E-02                  |                           |                           |+/-2.04E-02    |Jy       |1978ApJS...38..267O|uncertainty                   |2.28    microns    |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |9" aperture                             |Averaged new and previously published data                                                                                                                         
 242   |K                   |7.2E+00               |+/-0.04      |mag                 |1.31E+14 |7.92E-01    |2.97E-02                  |2.97E-02                  |                           |                           |+/-2.97E-02    |Jy       |1978ApJS...38..267O|uncertainty                   |2.28    microns    |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |18" aperture                            |Averaged new and previously published data                                                                                                                         
 246   |3.4 microns WISE AB |8.1E+00               |+/-0.10      |mag                 |8.93E+13 |2.06E+00    |1.90E-01                  |1.90E-01                  |                           |                           |+/-1.90E-01    |Jy       |2014ApJS..212...18B|uncertainty                   |33570   A          |Broad-band measurement                                                 |40.66969000 -0.01318000 (J2000)  |Flux in fixed aperture                                  |155"x180" aperture                      |From new raw data; Extinction-corrected for Milky Way                                                                                                              
 247   |3.4 microns WISE AB |8.1E+00               |+/-0.10      |mag                 |8.93E+13 |2.04E+00    |1.88E-01                  |1.88E-01                  |                           |                           |+/-1.88E-01    |Jy       |2014ApJS..212...18B|uncertainty                   |33570   A          |Broad-band measurement                                                 |40.66969000 -0.01318000 (J2000)  |Flux in fixed aperture                                  |155"x180" aperture                      |From new raw data                                                                                                                                                  
 248   |3.4 microns         |2.9E+00               |+/-0.3       |Jy                  |8.82E+13 |2.90E+00    |3.00E-01                  |3.00E-01                  |                           |                           |+/-3.00E-01    |Jy       |1970ApJ...159L.165K|no uncertainty reported       |3.4 microns        |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |                                        |From new raw data                                                                                                                                                  
 249   |3.4 microns         |5.4E+00               |+/-0.10      |mag                 |8.82E+13 |1.97E+00    |1.90E-01                  |1.90E-01                  |                           |                           |+/-1.90E-01    |Jy       |1974MNRAS.169..357P|uncertainty                   |3.4   microns      |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |10.0" aperture                          |From new raw data                                                                                                                                                  
 250   |3.4 microns         |5.3E+00               |+/-0.11      |mag                 |8.82E+13 |2.18E+00    |2.33E-01                  |2.33E-01                  |                           |                           |+/-2.33E-01    |Jy       |1974MNRAS.169..357P|uncertainty                   |3.4   microns      |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |32" aperture                            |From new raw data                                                                                                                                                  
 251   |3.4 microns         |5.2E+00               |+/-0.15      |mag                 |8.82E+13 |2.27E+00    |3.36E-01                  |3.36E-01                  |                           |                           |+/-3.36E-01    |Jy       |1974MNRAS.169..357P|uncertainty                   |3.4   microns      |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |22" aperture                            |From new raw data                                                                                                                                                  
 252   |3.4 microns         |5.4E+00               |             |mag                 |8.82E+13 |1.97E+00    |                          |                          |                           |                           |               |Jy       |1974MNRAS.169..357P|no uncertainty reported       |3.4   microns      |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |13.5" aperture                          |Averaged new and previously published data                                                                                                                         
 253   |3.4 microns         |5.3E+00               |             |mag                 |8.82E+13 |2.18E+00    |                          |                          |                           |                           |               |Jy       |1974MNRAS.169..357P|no uncertainty reported       |3.4   microns      |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |15" aperture                            |Averaged new and previously published data                                                                                                                         
 254   |3.4 microns         |5.3E+00               |+/-0.15      |mag                 |8.82E+13 |2.10E+00    |3.12E-01                  |3.12E-01                  |                           |                           |+/-3.12E-01    |Jy       |1974MNRAS.169..357P|uncertainty                   |3.4   microns      |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |20" aperture                            |From new raw data                                                                                                                                                  
 255   |3.5 microns         |1.7E+00               |+/-0.2       |Jy                  |8.57E+13 |1.70E+00    |2.00E-01                  |2.00E-01                  |                           |                           |+/-2.00E-01    |Jy       |1972ApJ...176L..95R|1 sigma                       |3.5 microns        |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |6" aperture                             |From new raw data                                                                                                                                                  
 256   |L                   |5.4E+00               |+/-0.07      |mag                 |8.57E+13 |1.88E+00    |1.26E-01                  |1.26E-01                  |                           |                           |+/-1.26E-01    |Jy       |1978ApJS...38..267O|uncertainty                   |3.5     microns    |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |18" aperture                            |Averaged new and previously published data                                                                                                                         
 257   |3.5 microns         |5.5E+00               |+/-0.1       |mag                 |8.57E+13 |1.85E+00    |1.78E-01                  |1.78E-01                  |                           |                           |+/-1.78E-01    |Jy       |1976ApJ...205...44S|uncertainty                   |3.5     microns    |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |8.4" aperture                           |Averaged new and previously published data                                                                                                                         
 258   |L                   |5.4E+00               |+/-0.07      |mag                 |8.57E+13 |1.88E+00    |1.26E-01                  |1.26E-01                  |                           |                           |+/-1.26E-01    |Jy       |1978ApJS...38..267O|uncertainty                   |3.5     microns    |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |9" aperture                             |Averaged new and previously published data                                                                                                                         
 259   |L (RGO)             |5.5E+00               |+/-0.03      |mag                 |8.57E+13 |1.72E+00    |4.82E-02                  |4.82E-02                  |                           |                           |+/-4.82E-02    |Jy       |1981MNRAS.197.1067G|uncertainty                   |3.5     microns    |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |12" aperture                            |From new raw data                                                                                                                                                  
 260   |L (Johnson)         |5.3E+00               |+/-0.1       |mag                 |8.47E+13 |2.19E+00    |2.11E-01                  |2.11E-01                  |                           |                           |+/-2.11E-01    |Jy       |1967ApJ...147..394P|uncertainty                   |3.54 microns       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |15" aperture                            |From new raw data                                                                                                                                                  
 261   |3.6 microns (IRAC)  |3.8E+00               |             |Jy                  |8.44E+13 |3.80E+00    |                          |                          |                           |                           |               |Jy       |2007AJ....134.2086H|no uncertainty reported       |3.550 microns      |Broad-band measurement                                                 |                                 |Total flux                                              |                                        |From new raw data                                                                                                                                                  
 262   |3.6 microns         |1.9E+00               |+/-10  %     |Jy                  |8.33E+13 |1.92E+00    |1.93E-01                  |1.93E-01                  |                           |                           |+/-1.93E-01    |Jy       |1978ApJ...226..550R|uncertainty                   |3.6     microns    |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |8.5" aperture                           |From new raw data                                                                                                                                                  
 265   |L (VLT)             |1.5E+00               |             |Jy                  |7.90E+13 |1.50E+00    |                          |                          |                           |                           |               |Jy       |2008A&A...485...33H|no uncertainty reported       |3.8 microns        |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |Nuclear flux                            |Averaged from previously published data                                                                                                                            
 266   |L' (VLT/NACO)       |8.8E+00               |             |mag                 |7.89E+13 |7.61E-02    |                          |                          |                           |                           |               |Jy       |2006A&A...446..813G|no uncertainty reported       |3.80   microns     |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |Nuclear; aperture radius = 0.08"        |From reprocessed raw data; derived from a flux in a differentband and a color                                                                                      
 267   |L' (VLT/NACO)       |6.6E+00               |             |mag                 |7.89E+13 |5.77E-01    |                          |                          |                           |                           |               |Jy       |2006A&A...446..813G|no uncertainty reported       |3.80   microns     |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |Nuclear; aperture radius = 0.27"        |From reprocessed raw data; derived from a flux in a differentband and a color                                                                                      
 268   |L' (VLT/NACO)       |7.7E+00               |             |mag                 |7.89E+13 |2.10E-01    |                          |                          |                           |                           |               |Jy       |2006A&A...446..813G|no uncertainty reported       |3.80   microns     |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |Nuclear; aperture radius = 0.13"        |From reprocessed raw data; derived from a flux in a differentband and a color                                                                                      
 271   |M (VLT)             |2.5E+00               |             |Jy                  |6.70E+13 |2.50E+00    |                          |                          |                           |                           |               |Jy       |2008A&A...485...33H|no uncertainty reported       |4.5  microns       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |Nuclear flux                            |From new raw data                                                                                                                                                  
 272   |4.5 microns (IRAC)  |5.1E+00               |             |Jy                  |6.67E+13 |5.10E+00    |                          |                          |                           |                           |               |Jy       |2007AJ....134.2086H|no uncertainty reported       |4.493 microns      |Broad-band measurement                                                 |                                 |Total flux                                              |                                        |From new raw data                                                                                                                                                  
 273   |4.5 microns (ISOCAM)|6.9E+03               |+/-340       |milliJy             |6.66E+13 |6.86E+00    |3.40E-01                  |3.40E-01                  |                           |                           |+/-3.40E-01    |Jy       |2004A&A...421..129S|1 sigma                       |4.5   microns      |Broad-band measurement                                                 |                                 |From multi-aperture data                                |                                        |From reprocessed raw data                                                                                                                                          
 275   |4.6 microns WISE AB |7.7E+00               |+/-0.10      |mag                 |6.51E+13 |2.98E+00    |2.74E-01                  |2.74E-01                  |                           |                           |+/-2.74E-01    |Jy       |2014ApJS..212...18B|uncertainty                   |46060   A          |Broad-band measurement                                                 |40.66969000 -0.01318000 (J2000)  |Flux in fixed aperture                                  |155"x180" aperture                      |From new raw data                                                                                                                                                  
 276   |4.6 microns WISE AB |7.7E+00               |+/-0.10      |mag                 |6.51E+13 |3.00E+00    |2.76E-01                  |2.76E-01                  |                           |                           |+/-2.76E-01    |Jy       |2014ApJS..212...18B|uncertainty                   |46060   A          |Broad-band measurement                                                 |40.66969000 -0.01318000 (J2000)  |Flux in fixed aperture                                  |155"x180" aperture                      |From new raw data; Extinction-corrected for Milky Way                                                                                                              
 278   |M' (VLT/NACO)       |5.6E+00               |             |mag                 |6.27E+13 |9.78E-01    |                          |                          |                           |                           |               |Jy       |2006A&A...446..813G|no uncertainty reported       |4.78   microns     |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |Nuclear; aperture radius = 0.13"        |From reprocessed raw data; derived from a flux in a differentband and a color                                                                                      
 279   |M' (VLT/NACO)       |4.9E+00               |             |mag                 |6.27E+13 |1.86E+00    |                          |                          |                           |                           |               |Jy       |2006A&A...446..813G|no uncertainty reported       |4.78   microns     |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |Nuclear; aperture radius = 0.27"        |From reprocessed raw data; derived from a flux in a differentband and a color                                                                                      
 280   |M' (VLT/NACO)       |6.6E+00               |             |mag                 |6.27E+13 |3.89E-01    |                          |                          |                           |                           |               |Jy       |2006A&A...446..813G|no uncertainty reported       |4.78   microns     |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |Nuclear; aperture radius = 0.08"        |From reprocessed raw data; derived from a flux in a differentband and a color                                                                                      
 281   |5.0 microns         |7.2E+00               |+/-0.3       |Jy                  |6.00E+13 |7.20E+00    |3.00E-01                  |3.00E-01                  |                           |                           |+/-3.00E-01    |Jy       |1970ApJ...159L.165K|no uncertainty reported       |5.0 microns        |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |Low quality data                        |From new raw data                                                                                                                                                  
 282   |5.0 microns         |3.2E+00               |+/-0.2       |Jy                  |6.00E+13 |3.20E+00    |2.00E-01                  |2.00E-01                  |                           |                           |+/-2.00E-01    |Jy       |1972ApJ...176L..95R|1 sigma                       |5.0 microns        |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |6" aperture                             |From new raw data                                                                                                                                                  
 283   |5.8 microns (IRAC)  |1.3E+01               |             |Jy                  |5.23E+13 |1.30E+01    |                          |                          |                           |                           |               |Jy       |2007AJ....134.2086H|no uncertainty reported       |5.731 microns      |Broad-band measurement                                                 |                                 |Total flux                                              |                                        |From new raw data                                                                                                                                                  
 284   |6 microns (ISO)     |1.1E+01               |             |Jy                  |5.00E+13 |1.12E+01    |                          |                          |                           |                           |               |Jy       |2004A&A...418..465L|no uncertainty reported       |6   microns        |Broad-band measurement                                                 |                                 |Flux integrated from map                                |                                        |From reprocessed raw data                                                                                                                                          
 285   |6.8 microns (ISOCAM)|1.4E+04               |+/-700       |milliJy             |4.41E+13 |1.40E+01    |7.00E-01                  |7.00E-01                  |                           |                           |+/-7.00E-01    |Jy       |2004A&A...421..129S|1 sigma                       |6.8   microns      |Broad-band measurement                                                 |                                 |From multi-aperture data                                |                                        |From reprocessed raw data                                                                                                                                          
 286   |8.0 microns (IRAC)  |2.3E+01               |             |Jy                  |3.81E+13 |2.30E+01    |                          |                          |                           |                           |               |Jy       |2007AJ....134.2086H|no uncertainty reported       |7.872 microns      |Broad-band measurement                                                 |                                 |Total flux                                              |                                        |From new raw data                                                                                                                                                  
 287   |8.6 microns TIMMI2  |1.5E+01               |+/-10  %     |Jy                  |3.49E+13 |1.48E+01    |1.48E+00                  |1.48E+00                  |                           |                           |+/-1.48E+00    |Jy       |2004A&A...414..123S|uncertainty                   |8.6   microns      |Broad-band measurement                                                 |                                 |From multi-aperture data                                |                                        |From new raw data                                                                                                                                                  
 288   |PAH1 (VLT)          |1.9E+04               |+/-657.0     |milliJy             |3.49E+13 |1.85E+01    |6.57E-01                  |6.57E-01                  |                           |                           |+/-6.57E-01    |Jy       |2014MNRAS.439.1648A|uncertainty                   |8.59   microns     |Broad-band measurement                                                 |040.669583 -00.013333 (J2000)    |Flux in fixed aperture                                  |Nuclear flux                            |From reprocessed raw data                                                                                                                                          
 289   |8.99 microns (VLT)  |6.8E+00               |+/-0.2       |Jy                  |3.33E+13 |6.80E+00    |2.00E-01                  |2.00E-01                  |                           |                           |+/-2.00E-01    |Jy       |2008A&A...481..305P|estimated error               |8.99 microns       |Broad-band measurement                                                 |                                 |From fitting to map                                     |Slit at -15deg                          |From new raw data                                                                                                                                                  
 290   |8.99 microns (VLT)  |7.8E+00               |+/-0.4       |Jy                  |3.33E+13 |7.80E+00    |4.00E-01                  |4.00E-01                  |                           |                           |+/-4.00E-01    |Jy       |2008A&A...481..305P|estimated error               |8.99 microns       |Broad-band measurement                                                 |                                 |From fitting to map                                     |Slit at 90deg                           |From new raw data                                                                                                                                                  
 291   |ARIII (VLT)         |1.8E+04               |+/-469.0     |milliJy             |3.33E+13 |1.78E+01    |4.69E-01                  |4.69E-01                  |                           |                           |+/-4.69E-01    |Jy       |2014MNRAS.439.1648A|uncertainty                   |8.99   microns     |Broad-band measurement                                                 |040.669583 -00.013333 (J2000)    |Flux in fixed aperture                                  |Nuclear flux                            |From reprocessed raw data                                                                                                                                          
 292   |10 microns          |2.5E+01               |+/-3         |Jy                  |3.00E+13 |2.50E+01    |3.00E+00                  |3.00E+00                  |                           |                           |+/-3.00E+00    |Jy       |1972ApJ...177L.115R|uncertainty                   |10 microns         |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |6" aperture;Low quality data            |From new raw data                                                                                                                                                  
 293   |10 microns          |2.5E+01               |             |Jy                  |3.00E+13 |2.50E+01    |                          |                          |                           |                           |               |Jy       |1978ApJ...220L..37R|no uncertainty reported       |10      microns    |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |5.7" aperture                           |From new raw data                                                                                                                                                  
 294   |10.2 microns        |3.1E+01               |+/-0.2       |Jy                  |2.94E+13 |3.06E+01    |2.00E-01                  |2.00E-01                  |                           |                           |+/-2.00E-01    |Jy       |1970ApJ...159L.165K|no uncertainty reported       |10.2 microns       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |Low quality data                        |From new raw data                                                                                                                                                  
 295   |10.4 microns TIMMI2 |1.8E+01               |+/-10  %     |Jy                  |2.88E+13 |1.76E+01    |1.76E+00                  |1.76E+00                  |                           |                           |+/-1.76E+00    |Jy       |2004A&A...414..123S|uncertainty                   |10.4   microns     |Broad-band measurement                                                 |                                 |From multi-aperture data                                |                                        |From new raw data                                                                                                                                                  
 296   |10.5 microns        |2.5E+01               |             |Jy                  |2.86E+13 |2.50E+01    |                          |                          |                           |                           |               |Jy       |1972ApJ...176L..95R|no uncertainty reported       |10.5 microns       |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |6" aperture                             |From new raw data                                                                                                                                                  
 300   |10.51 microns (VLT) |8.3E+00               |+/-0.2       |Jy                  |2.85E+13 |8.30E+00    |2.00E-01                  |2.00E-01                  |                           |                           |+/-2.00E-01    |Jy       |2008A&A...481..305P|estimated error               |10.51 microns      |Broad-band measurement                                                 |                                 |From fitting to map                                     |Slit at -15deg                          |From new raw data                                                                                                                                                  
 301   |10.51 microns (VLT) |1.0E+01               |+/-0.3       |Jy                  |2.85E+13 |1.02E+01    |3.00E-01                  |3.00E-01                  |                           |                           |+/-3.00E-01    |Jy       |2008A&A...481..305P|estimated error               |10.51 microns      |Broad-band measurement                                                 |                                 |From fitting to map                                     |Slit at 90deg                           |From new raw data                                                                                                                                                  
 303   |10.6 microns        |1.8E+01               |+/-10  %     |Jy                  |2.83E+13 |1.80E+01    |1.80E+00                  |1.80E+00                  |                           |                           |+/-1.80E+00    |Jy       |1978ApJ...226..550R|uncertainty                   |10.6     microns   |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |5.7" aperture                           |From new raw data                                                                                                                                                  
 304   |10.6 microns        |1.8E+01               |             |Jy                  |2.83E+13 |1.80E+01    |                          |                          |                           |                           |               |Jy       |1979ApJ...229..111L|no uncertainty reported       |10.6     microns   |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |8.5" aperture                           |From new raw data                                                                                                                                                  
 305   |N (Johnson)         |9.6E-01               |+/-0.16      |mag                 |2.83E+13 |1.49E+01    |2.36E+00                  |2.36E+00                  |                           |                           |+/-2.36E+00    |Jy       |1983ApJ...275..477M|uncertainty                   |10.6     microns   |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |9" aperture                             |From new raw data                                                                                                                                                  
 306   |10.8 microns MIRLIN |2.6E+04               |+/-3200      |milliJy             |2.78E+13 |2.56E+01    |3.20E+00                  |3.20E+00                  |                           |                           |+/-3.20E+00    |Jy       |2004ApJ...605..156G|statistical error             |10.8   microns     |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |1.5" diam aperture                      |From new raw data                                                                                                                                                  
 307   |SIV_2 (VLT)         |2.7E+04               |+/-773.3     |milliJy             |2.78E+13 |2.68E+01    |7.73E-01                  |7.73E-01                  |                           |                           |+/-7.73E-01    |Jy       |2014MNRAS.439.1648A|uncertainty                   |10.77   microns    |Broad-band measurement                                                 |040.669583 -00.013333 (J2000)    |Flux in fixed aperture                                  |Nuclear flux                            |From reprocessed raw data                                                                                                                                          
 308   |PAH2 (VLT)          |2.9E+04               |+/-653.8     |milliJy             |2.66E+13 |2.92E+01    |6.54E-01                  |6.54E-01                  |                           |                           |+/-6.54E-01    |Jy       |2014MNRAS.439.1648A|uncertainty                   |11.25   microns    |Broad-band measurement                                                 |040.669583 -00.013333 (J2000)    |Flux in fixed aperture                                  |Nuclear flux                            |From reprocessed raw data                                                                                                                                          
 311   |SIC (VLT)           |3.2E+04               |+/-1789.8    |milliJy             |2.53E+13 |3.18E+01    |1.79E+00                  |1.79E+00                  |                           |                           |+/-1.79E+00    |Jy       |2014MNRAS.439.1648A|uncertainty                   |11.85   microns    |Broad-band measurement                                                 |040.669583 -00.013333 (J2000)    |Flux in fixed aperture                                  |Nuclear flux                            |From reprocessed raw data                                                                                                                                          
 312   |12 microns (IRAS)   |4.0E+01               |+/-0.076     |Jy                  |2.50E+13 |3.98E+01    |7.60E-02                  |7.60E-02                  |                           |                           |+/-7.60E-02    |Jy       |2003AJ....126.1607S|1 sigma                       |12   microns       |Broad-band measurement                                                 |02 42 41.4 -00 00 45 (J2000)     |Total flux                                              |Size, Method, Flag codes: MI;see paper  |From reprocessed raw data                                                                                                                                          
 313   |12 microns (VLTI)   |1.7E+01               |             |Jy                  |2.50E+13 |1.65E+01    |                          |                          |                           |                           |               |Jy       |2009A&A...502...67T|no uncertainty reported       |12 microns         |Broad-band measurement                                                 |02 42 40.70 -00 00 48.0 (J2000)  |Total flux                                              |                                        |From new raw data                                                                                                                                                  
 314   |12 microns (IRAS)   |3.9E+04               |+/-15  %     |milliJy             |2.50E+13 |3.87E+01    |5.80E+00                  |5.80E+00                  |                           |                           |+/-5.80E+00    |Jy       |1988AJ.....95...26G|typical accuracy              |12         microns |Broad-band measurement                                                 |                                 |Integrated from scans                                   |From pointed observations               |From new raw data                                                                                                                                                  
 315   |12 microns (IRAS)   |3.6E+01               |+/-0.064     |Jy                  |2.50E+13 |3.61E+01    |6.40E-02                  |6.40E-02                  |                           |                           |+/-6.40E-02    |Jy       |1989AJ.....98..766S|rms noise                     |12         microns |Broad-band measurement                                                 |024007.2 -001330 (B1950)         |Integrated from scans                                   |Unresolved with 0.77' beam              |From reprocessed raw data                                                                                                                                          
 316   |12 microns (IRAS)   |4.0E+01               |+/-5   %     |Jy                  |2.50E+13 |3.97E+01    |1.99E+00                  |1.99E+00                  |                           |                           |+/-1.99E+00    |Jy       |1990IRASF.C...0000M|uncertainty                   |12        microns  |Broad-band measurement                                                 |024007.7 -001329 (B1950)         |Flux in fixed aperture                                  |IRAS quality flag = 3                   |From new raw data                                                                                                                                                  
 317   |NEII_1 (VLT)        |3.2E+04               |+/-822.7     |milliJy             |2.44E+13 |3.18E+01    |8.23E-01                  |8.23E-01                  |                           |                           |+/-8.23E-01    |Jy       |2014MNRAS.439.1648A|uncertainty                   |12.27   microns    |Broad-band measurement                                                 |040.669583 -00.013333 (J2000)    |Flux in fixed aperture                                  |Nuclear flux                            |From reprocessed raw data                                                                                                                                          
 319   |12.81 microns (VLT) |1.3E+01               |+/-0.5       |Jy                  |2.34E+13 |1.28E+01    |5.00E-01                  |5.00E-01                  |                           |                           |+/-5.00E-01    |Jy       |2008A&A...481..305P|estimated error               |12.81 microns      |Broad-band measurement                                                 |                                 |From fitting to map                                     |Slit at -15deg                          |From new raw data                                                                                                                                                  
 320   |12.81 microns (VLT) |1.7E+01               |+/-1.2       |Jy                  |2.34E+13 |1.72E+01    |1.20E+00                  |1.20E+00                  |                           |                           |+/-1.20E+00    |Jy       |2008A&A...481..305P|estimated error               |12.81 microns      |Broad-band measurement                                                 |                                 |From fitting to map                                     |Slit at 90deg                           |From new raw data                                                                                                                                                  
 327   |NEII (VLT)          |3.7E+04               |+/-1317.6    |milliJy             |2.34E+13 |3.65E+01    |1.32E+00                  |1.32E+00                  |                           |                           |+/-1.32E+00    |Jy       |2014MNRAS.439.1648A|uncertainty                   |12.81   microns    |Broad-band measurement                                                 |040.669583 -00.013333 (J2000)    |Flux in fixed aperture                                  |Nuclear flux                            |From reprocessed raw data                                                                                                                                          
 328   |NEII_2 (VLT)        |3.5E+04               |+/-1403.4    |milliJy             |2.30E+13 |3.52E+01    |1.40E+00                  |1.40E+00                  |                           |                           |+/-1.40E+00    |Jy       |2014MNRAS.439.1648A|uncertainty                   |13.04   microns    |Broad-band measurement                                                 |040.669583 -00.013333 (J2000)    |Flux in fixed aperture                                  |Nuclear flux                            |From reprocessed raw data                                                                                                                                          
 335   |14.9 microns ISOCAM |5.1E+04               |+/-2540      |milliJy             |2.01E+13 |5.08E+01    |2.54E+00                  |2.54E+00                  |                           |                           |+/-2.54E+00    |Jy       |2004A&A...421..129S|1 sigma                       |14.9   microns     |Broad-band measurement                                                 |                                 |From multi-aperture data                                |                                        |From reprocessed raw data                                                                                                                                          
 341   |Q1 (VLT)            |5.8E+04               |+/-1243.6    |milliJy             |1.70E+13 |5.76E+01    |1.24E+00                  |1.24E+00                  |                           |                           |+/-1.24E+00    |Jy       |2014MNRAS.439.1648A|uncertainty                   |17.65   microns    |Broad-band measurement                                                 |040.669583 -00.013333 (J2000)    |Flux in fixed aperture                                  |Nuclear flux                            |From reprocessed raw data                                                                                                                                          
 343   |Q2 (VLT)            |6.7E+04               |+/-2030.0    |milliJy             |1.60E+13 |6.69E+01    |2.03E+00                  |2.03E+00                  |                           |                           |+/-2.03E+00    |Jy       |2014MNRAS.439.1648A|uncertainty                   |18.72   microns    |Broad-band measurement                                                 |040.669583 -00.013333 (J2000)    |Flux in fixed aperture                                  |Nuclear flux                            |From reprocessed raw data                                                                                                                                          
 344   |Q3 (VLT)            |5.7E+04               |+/-1662.9    |milliJy             |1.54E+13 |5.75E+01    |1.66E+00                  |1.66E+00                  |                           |                           |+/-1.66E+00    |Jy       |2014MNRAS.439.1648A|uncertainty                   |19.50   microns    |Broad-band measurement                                                 |040.669583 -00.013333 (J2000)    |Flux in fixed aperture                                  |Nuclear flux                            |From reprocessed raw data                                                                                                                                          
 345   |21 microns          |5.6E+01               |+/-4         |Jy                  |1.43E+13 |5.60E+01    |4.00E+00                  |4.00E+00                  |                           |                           |+/-4.00E+00    |Jy       |1972ApJ...176L..95R|1 sigma                       |21 microns         |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |6" aperture                             |From new raw data                                                                                                                                                  
 346   |21 microns          |6.6E+01               |             |Jy                  |1.43E+13 |6.60E+01    |                          |                          |                           |                           |               |Jy       |1979ApJ...229..111L|no uncertainty reported       |21       microns   |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |8.5" aperture                           |Recalibrated data                                                                                                                                                  
 347   |22 microns          |8.0E+01               |+/-5         |Jy                  |1.36E+13 |8.00E+01    |5.00E+00                  |5.00E+00                  |                           |                           |+/-5.00E+00    |Jy       |1970ApJ...159L.165K|no uncertainty reported       |22 microns         |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |                                        |From new raw data                                                                                                                                                  
 348   |22 microns WISE AB  |4.5E+00               |+/-0.10      |mag                 |1.35E+13 |5.62E+01    |5.18E+00                  |5.18E+00                  |                           |                           |+/-5.18E+00    |Jy       |2014ApJS..212...18B|uncertainty                   |221400   A         |Broad-band measurement                                                 |40.66969000 -0.01318000 (J2000)  |Flux in fixed aperture                                  |155"x180" aperture                      |From new raw data; Extinction-corrected for Milky Way                                                                                                              
 349   |22 microns WISE AB  |4.5E+00               |+/-0.10      |mag                 |1.35E+13 |5.62E+01    |5.17E+00                  |5.17E+00                  |                           |                           |+/-5.17E+00    |Jy       |2014ApJS..212...18B|uncertainty                   |221400   A         |Broad-band measurement                                                 |40.66969000 -0.01318000 (J2000)  |Flux in fixed aperture                                  |155"x180" aperture                      |From new raw data                                                                                                                                                  
 350   |24 microns (MIPS)   |8.0E+01               |             |Jy                  |1.27E+13 |8.00E+01    |                          |                          |                           |                           |               |Jy       |2007AJ....134.2086H|no uncertainty reported       |23.68 microns      |Broad-band measurement                                                 |                                 |Total flux                                              |                                        |From new raw data                                                                                                                                                  
 354   |25 microns (IRAS)   |8.8E+01               |+/-0.171     |Jy                  |1.20E+13 |8.76E+01    |1.71E-01                  |1.71E-01                  |                           |                           |+/-1.71E-01    |Jy       |2003AJ....126.1607S|1 sigma                       |25   microns       |Broad-band measurement                                                 |02 42 41.4 -00 00 45 (J2000)     |Total flux                                              |Size, Method, Flag codes: UT;see paper  |From reprocessed raw data                                                                                                                                          
 355   |25 microns (IRAS)   |8.7E+04               |+/-15  %     |milliJy             |1.20E+13 |8.74E+01    |1.31E+01                  |1.31E+01                  |                           |                           |+/-1.31E+01    |Jy       |1988AJ.....95...26G|typical accuracy              |25         microns |Broad-band measurement                                                 |                                 |Integrated from scans                                   |From pointed observations               |From new raw data                                                                                                                                                  
 356   |25 microns (IRAS)   |8.4E+01               |+/-0.191     |Jy                  |1.20E+13 |8.42E+01    |1.91E-01                  |1.91E-01                  |                           |                           |+/-1.91E-01    |Jy       |1989AJ.....98..766S|rms noise                     |25         microns |Broad-band measurement                                                 |024007.2 -001330 (B1950)         |Integrated from scans                                   |Unresolved with 0.78' beam              |From reprocessed raw data                                                                                                                                          
 357   |25 microns (IRAS)   |8.5E+01               |+/-6   %     |Jy                  |1.20E+13 |8.50E+01    |2.38E+00                  |2.38E+00                  |                           |                           |+/-2.38E+00    |Jy       |1990IRASF.C...0000M|uncertainty                   |25        microns  |Broad-band measurement                                                 |024007.7 -001329 (B1950)         |Flux in fixed aperture                                  |IRAS quality flag = 3                   |From new raw data                                                                                                                                                  
 374   |60 microns (IRAS)   |1.8E+05               |+/-15  %     |milliJy             |5.00E+12 |1.75E+02    |2.62E+01                  |2.62E+01                  |                           |                           |+/-2.62E+01    |Jy       |1988AJ.....95...26G|typical accuracy              |60         microns |Broad-band measurement                                                 |                                 |Integrated from scans                                   |From pointed observations               |From new raw data                                                                                                                                                  
 375   |60 microns (IRAS)   |2.0E+02               |+/-0.108     |Jy                  |5.00E+12 |1.96E+02    |1.08E-01                  |1.08E-01                  |                           |                           |+/-1.08E-01    |Jy       |2003AJ....126.1607S|1 sigma                       |60   microns       |Broad-band measurement                                                 |02 42 41.4 -00 00 45 (J2000)     |Total flux                                              |Size, Method, Flag codes: MI;see paper  |From reprocessed raw data                                                                                                                                          
 376   |60 microns (ISO)    |2.1E+02               |+/-20  %     |Jy                  |5.00E+12 |2.06E+02    |4.13E+01                  |4.13E+01                  |                           |                           |+/-4.13E+01    |Jy       |2001A&A...375..566N|uncertainty                   |60   microns       |Broad-band measurement                                                 |                                 |Modelled datum                                          |                                        |From new raw data                                                                                                                                                  
 377   |60 microns (IRAS)   |1.8E+02               |+/-0.103     |Jy                  |5.00E+12 |1.82E+02    |1.03E-01                  |1.03E-01                  |                           |                           |+/-1.03E-01    |Jy       |1989AJ.....98..766S|rms noise                     |60         microns |Broad-band measurement                                                 |024007.2 -001330 (B1950)         |Integrated from scans                                   |Unresolved with 1.44' beam              |From reprocessed raw data                                                                                                                                          
 378   |60 microns (IRAS)   |1.8E+02               |+/-5   %     |Jy                  |5.00E+12 |1.76E+02    |8.81E+00                  |8.81E+00                  |                           |                           |+/-8.81E+00    |Jy       |1990IRASF.C...0000M|uncertainty                   |60        microns  |Broad-band measurement                                                 |024007.7 -001329 (B1950)         |Flux in fixed aperture                                  |IRAS quality flag = 3                   |From new raw data                                                                                                                                                  
 381   |70 microns (MIPS)   |1.8E+02               |             |Jy                  |4.20E+12 |1.80E+02    |                          |                          |                           |                           |               |Jy       |2007AJ....134.2086H|no uncertainty reported       |71.42 microns      |Broad-band measurement                                                 |                                 |Total flux                                              |                                        |From new raw data                                                                                                                                                  
 383   |88 microns          |3.3E+02               |+/-74        |Jy                  |3.41E+12 |3.30E+02    |7.40E+01                  |7.40E+01                  |                           |                           |+/-7.40E+01    |Jy       |1977ApJ...216..698H|estimated error               |88        microns  |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |Beam diameter 45 arcsec                 |From new raw data                                                                                                                                                  
 384   |100 microns (IRAS)  |2.8E+05               |+/-15  %     |milliJy             |3.00E+12 |2.77E+02    |4.16E+01                  |4.16E+01                  |                           |                           |+/-4.16E+01    |Jy       |1988AJ.....95...26G|typical accuracy              |100        microns |Broad-band measurement                                                 |                                 |Integrated from scans                                   |From pointed observations               |From new raw data                                                                                                                                                  
 385   |100 microns (IRAS)  |2.6E+02               |+/-0.228     |Jy                  |3.00E+12 |2.57E+02    |2.28E-01                  |2.28E-01                  |                           |                           |+/-2.28E-01    |Jy       |2003AJ....126.1607S|1 sigma                       |100   microns      |Broad-band measurement                                                 |02 42 41.4 -00 00 45 (J2000)     |Total flux                                              |Size, Method, Flag codes: MI;see paper  |From reprocessed raw data                                                                                                                                          
 386   |100 microns (IRAS)  |2.2E+02               |+/-4   %     |Jy                  |3.00E+12 |2.24E+02    |8.96E+00                  |8.96E+00                  |                           |                           |+/-8.96E+00    |Jy       |1990IRASF.C...0000M|uncertainty                   |100       microns  |Broad-band measurement                                                 |024007.7 -001329 (B1950)         |Flux in fixed aperture                                  |IRAS quality flag = 2                   |From new raw data                                                                                                                                                  
 387   |100 microns (IRAS)  |2.4E+02               |+/-0.218     |Jy                  |3.00E+12 |2.36E+02    |2.18E-01                  |2.18E-01                  |                           |                           |+/-2.18E-01    |Jy       |1989AJ.....98..766S|rms noise                     |100        microns |Broad-band measurement                                                 |024007.2 -001330 (B1950)         |Integrated from scans                                   |Unresolved with 2.94' beam              |From reprocessed raw data                                                                                                                                          
 389   |134 microns         |2.7E+02               |+/-92        |Jy                  |2.24E+12 |2.72E+02    |9.20E+01                  |9.20E+01                  |                           |                           |+/-9.20E+01    |Jy       |1977ApJ...216..698H|estimated error               |134       microns  |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |Beam diameter 45 arcsec                 |From new raw data                                                                                                                                                  
 394   |170 microns (ISO)   |                      |>99.1        |Jy                  |1.76E+12 |            |                          |                          |                           |99.10000000                |>9.91E+01      |Jy       |2004A&A...422...39S|no uncertainty reported       |170      microns   |Broad-band measurement                                                 |02 42 40.7 -00 00 48 (J2000)     |Integrated from scans                                   |                                        |Averaged from previously published data                                                                                                                            
 395   |170 microns (ISO)   |3.9E+02               |+/-15  %     |Jy                  |1.76E+12 |3.89E+02    |5.84E+01                  |5.84E+01                  |                           |                           |+/-5.84E+01    |Jy       |2004A&A...422...39S|uncertainty                   |170      microns   |Broad-band measurement                                                 |02 42 40.54 -00 00 50.1 (J2000)  |Integrated from scans                                   |                                        |Averaged from previously published data                                                                                                                            
 396   |350 microns         |3.3E+01               |+/-0.82      |Jy                  |8.57E+11 |3.25E+01    |8.20E-01                  |8.20E-01                  |                           |                           |+/-8.20E-01    |Jy       |1999CIT...T00R....B|1 sigma                       |350        microns |Broad-band measurement                                                 |                                 |Flux integrated from map                                |                                        |From new raw data                                                                                                                                                  
 397   |390 microns         |3.0E+01               |+/-10        |Jy                  |7.69E+11 |3.00E+01    |1.00E+01                  |1.00E+01                  |                           |                           |+/-1.00E+01    |Jy       |1977ApJ...216..698H|based on count statistics only|390       microns  |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |Beam diameter 76 arcsec                 |From new raw data                                                                                                                                                  
 398   |390 microns         |3.3E+01               |+/-7         |Jy                  |7.69E+11 |3.30E+01    |7.00E+00                  |7.00E+00                  |                           |                           |+/-7.00E+00    |Jy       |1977ApJ...216..698H|based on count statistics only|390       microns  |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |Beam diameter 75 arcsec                 |From new raw data                                                                                                                                                  
 399   |540 microns         |                      |<7           |Jy                  |5.55E+11 |            |                          |                          |7.00000000                 |                           |<7.00E+00      |Jy       |1977ApJ...216..698H|2 sigma                       |540       microns  |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |Beam diameter 83 arcsec                 |From new raw data                                                                                                                                                  
 400   |810 microns (SMA)   |4.1E+01               |+/-11        |milliJy             |3.70E+11 |4.10E-02    |1.10E-02                  |1.10E-02                  |                           |                           |+/-1.10E-02    |Jy       |2011ApJ...736...37K|statistical error             |810 microns        |Broad-band measurement                                                 |02 42 40.70 -00 00 47.9 (J2000)  |From fitting to map                                     |Beam = 2.1" x 2.0"; PA = 80 deg         |From new raw data                                                                                                                                                  
 403   |850 microns (SMA)   |3.0E+01               |+/-5         |milliJy             |3.53E+11 |3.00E-02    |5.00E-03                  |5.00E-03                  |                           |                           |+/-5.00E-03    |Jy       |2011ApJ...736...37K|statistical error             |850 microns        |Broad-band measurement                                                 |02 42 40.70 -00 00 47.9 (J2000)  |From fitting to map                                     |Beam=0.6"x0.5";PA=30deg; unif. weighting|From new raw data                                                                                                                                                  
 404   |850 microns (SMA)   |5.0E+01               |+/-7         |milliJy             |3.53E+11 |5.00E-02    |7.00E-03                  |7.00E-03                  |                           |                           |+/-7.00E-03    |Jy       |2011ApJ...736...37K|statistical error             |850 microns        |Broad-band measurement                                                 |02 42 40.70 -00 00 47.9 (J2000)  |From fitting to map                                     |Beam=1.0"x0.8";PA=30deg; nat. weighting |From new raw data                                                                                                                                                  
 406   |1 mm (IRAM)         |2.2E+01               |+/-0.8       |milliJy             |3.00E+11 |2.20E-02    |8.00E-04                  |8.00E-04                  |                           |                           |+/-8.00E-04    |Jy       |2006A&A...446..113K|uncertainty                   |1   mm             |Broad-band measurement                                                 |                                 |Flux integrated from map                                |Core flux                               |From new raw data                                                                                                                                                  
 407   |1.0 mm (SMA)        |1.3E+01               |+/-2         |milliJy             |3.00E+11 |1.30E-02    |2.00E-03                  |2.00E-03                  |                           |                           |+/-2.00E-03    |Jy       |2011ApJ...736...37K|statistical error             |1.0 mm             |Broad-band measurement                                                 |02 42 40.70 -00 00 47.9 (J2000)  |From fitting to map                                     |Beam=0.5"x0.4";PA=30deg; unif. weighting|From new raw data                                                                                                                                                  
 408   |1.0 mm (SMA)        |2.4E+01               |+/-3         |milliJy             |3.00E+11 |2.40E-02    |3.00E-03                  |3.00E-03                  |                           |                           |+/-3.00E-03    |Jy       |2011ApJ...736...37K|statistical error             |1.0 mm             |Broad-band measurement                                                 |02 42 40.70 -00 00 47.9 (J2000)  |From fitting to map                                     |Beam=1.0"x0.8";PA=30deg; nat. weighting |From new raw data                                                                                                                                                  
 411   |1.3 mm (PdBI)       |2.2E+01               |+/-2         |milliJy             |2.31E+11 |2.20E-02    |2.00E-03                  |2.00E-03                  |                           |                           |+/-2.00E-03    |Jy       |2011ApJ...736...37K|statistical error             |1.3 mm             |Broad-band measurement                                                 |02 42 40.70 -00 00 47.9 (J2000)  |From fitting to map                                     |Beam = 1.0" x 0.8"; PA = 30 deg         |From new raw data                                                                                                                                                  
 413   |1.3 mm (NRAO)       |1.7E-01               |+/-0.03      |Jy                  |2.31E+11 |1.70E-01    |3.00E-02                  |3.00E-02                  |                           |                           |+/-3.00E-02    |Jy       |1987ApJ...318..645T|uncertainty                   |1.3 mm             |Broad-band measurement                                                 |02406.5 -001332 (B1950)          |Not reported in paper                                   |Beam size = 33"                         |From new raw data                                                                                                                                                  
 414   |1.4 mm (NIKA)       |1.4E+02               |+/-25        |milliJy             |2.20E+11 |1.42E-01    |2.50E-02                  |2.50E-02                  |                           |                           |+/-2.50E-02    |Jy       |2011ApJS..194...24M|uncertainty                   |1.4  mm            |Broad-band measurement                                                 |                                 |Flux integrated from map                                |Central flux                            |From new raw data                                                                                                                                                  
 417   |1.4 mm (SMA)        |2.8E+01               |+/-3         |milliJy             |2.14E+11 |2.80E-02    |3.00E-03                  |3.00E-03                  |                           |                           |+/-3.00E-03    |Jy       |2011ApJ...736...37K|statistical error             |1.4 mm             |Broad-band measurement                                                 |02 42 40.70 -00 00 47.9 (J2000)  |From fitting to map                                     |Beam = 1.0" x 0.8"; PA = 30 deg         |From new raw data                                                                                                                                                  
 418   |2 mm (NIKA)         |6.6E+01               |+/-3         |milliJy             |1.50E+11 |6.60E-02    |3.00E-03                  |3.00E-03                  |                           |                           |+/-3.00E-03    |Jy       |2011ApJS..194...24M|uncertainty                   |2    mm            |Broad-band measurement                                                 |                                 |Flux integrated from map                                |Central flux                            |From new raw data                                                                                                                                                  
 421   |3 mm (IRAM)         |3.6E+01               |+/-0.4       |milliJy             |9.99E+10 |3.60E-02    |4.00E-04                  |4.00E-04                  |                           |                           |+/-4.00E-04    |Jy       |2006A&A...446..113K|uncertainty                   |3   mm             |Broad-band measurement                                                 |                                 |Flux integrated from map                                |Core flux                               |From new raw data                                                                                                                                                  
 426   |43.34 GHz (VLA)     |1.8E+02               |+/-5.3       |milliJy             |4.33E+10 |1.75E-01    |5.30E-03                  |5.30E-03                  |                           |                           |+/-5.30E-03    |Jy       |2011ApJ...732...45S|rms uncertainty               |43.34 GHz          |Broad-band measurement                                                 |                                 |Total flux                                              |                                        |From new raw data                                                                                                                                                  
 427   |43.34 GHz (VLA)     |7.9E+01               |+/-2.1       |milliJy             |4.33E+10 |7.87E-02    |2.10E-03                  |2.10E-03                  |                           |                           |+/-2.10E-03    |Jy       |2011ApJ...732...45S|rms uncertainty               |43.34 GHz          |Broad-band measurement                                                 |                                 |Flux integrated from map                                |Core flux                               |From new raw data                                                                                                                                                  
 428   |43 GHz (VLA)        |2.1E+01               |+/-0.6       |milliJy             |4.30E+10 |2.12E-02    |6.00E-04                  |6.00E-04                  |                           |                           |+/-6.00E-04    |Jy       |2008A&A...477..517C|1 sigma                       |43   GHz           |Broad-band measurement                                                 |                                 |Flux integrated from map                                |Core flux                               |From new raw data                                                                                                                                                  
 429   |31 GHz (OVRO)       |3.2E+02               |+/-16.46     |milliJy             |3.10E+10 |3.17E-01    |1.65E-02                  |1.65E-02                  |                           |                           |+/-1.65E-02    |Jy       |2009ApJ...704.1433M|uncertainty                   |31 GHz             |Broad-band measurement                                                 |02 42 40.72 -00 00 47.7 (J2000)  |Flux integrated from map                                |                                        |From new raw data                                                                                                                                                  
 430   |25.1 GHz (GBT)      |3.7E-01               |             |Jy                  |2.51E+10 |3.70E-01    |                          |                          |                           |                           |               |Jy       |2011A&A...529A.154A|no uncertainty reported       |25.1 GHz           |Broad-band measurement                                                 |                                 |Flux integrated from map                                |                                        |From new raw data                                                                                                                                                  
 431   |23.4 GHz (GBT)      |3.3E-01               |             |Jy                  |2.34E+10 |3.30E-01    |                          |                          |                           |                           |               |Jy       |2011A&A...529A.154A|no uncertainty reported       |23.4 GHz           |Broad-band measurement                                                 |                                 |Flux integrated from map                                |                                        |From new raw data                                                                                                                                                  
 432   |23 GHz (WMAP)       |9.2E+02               |+/-158       |milliJy             |2.30E+10 |9.21E-01    |1.58E-01                  |1.58E-01                  |                           |                           |+/-1.58E-01    |Jy       |2009MNRAS.392..733M|uncertainty                   |23 GHz             |Broad-band measurement                                                 |040.5990 -00.0710 (J2000)        |Flux integrated from map                                |                                        |From new raw data                                                                                                                                                  
 433   |22.46 GHz (VLA)     |1.6E+02               |+/-2.0       |milliJy             |2.25E+10 |1.61E-01    |2.00E-03                  |2.00E-03                  |                           |                           |+/-2.00E-03    |Jy       |2011ApJ...732...45S|rms uncertainty               |22.46 GHz          |Broad-band measurement                                                 |                                 |Flux integrated from map                                |Core flux                               |From new raw data                                                                                                                                                  
 434   |22.46 GHz (VLA)     |3.2E+02               |+/-10.0      |milliJy             |2.25E+10 |3.20E-01    |1.00E-02                  |1.00E-02                  |                           |                           |+/-1.00E-02    |Jy       |2011ApJ...732...45S|rms uncertainty               |22.46 GHz          |Broad-band measurement                                                 |                                 |Total flux                                              |                                        |From new raw data                                                                                                                                                  
 435   |22 GHz (ATCA)       |3.4E-01               |+/-0.034     |Jy                  |2.20E+10 |3.42E-01    |3.40E-02                  |3.40E-02                  |                           |                           |+/-3.40E-02    |Jy       |2006A&A...445..465R|uncertainty                   |22   GHz           |Broad-band measurement                                                 |                                 |Modelled datum                                          |Resolved                                |From new raw data                                                                                                                                                  
 436   |20.0 GHz (OVRO)     |4.5E+02               |+/-34        |milliJy             |2.00E+10 |4.50E-01    |3.40E-02                  |3.40E-02                  |                           |                           |+/-3.40E-02    |Jy       |1987ApJ...313..651E|uncertainty                   |20.0   GHz         |Broad-band measurement                                                 |02 40 07.06 -00 13 30.3 (B1950)  |Flux integrated from map                                |                                        |From new raw data                                                                                                                                                  
 437   |20 GHz (ATCA)       |4.7E+02               |+/-17        |milliJy             |1.99E+10 |4.74E-01    |1.70E-02                  |1.70E-02                  |                           |                           |+/-1.70E-02    |Jy       |2010MNRAS.402.2403M|rms uncertainty               |19.904 GHz         |Broad-band measurement                                                 |02 42 40.72 -00 00 46.7 (J2000)  |Flux integrated from map                                |                                        |From new raw data                                                                                                                                                  
 438   |18.5 GHz (ATCA)     |4.3E-01               |+/-0.022     |Jy                  |1.85E+10 |4.32E-01    |2.20E-02                  |2.20E-02                  |                           |                           |+/-2.20E-02    |Jy       |2006A&A...445..465R|uncertainty                   |18.5   GHz         |Broad-band measurement                                                 |                                 |Modelled datum                                          |Resolved                                |From new raw data                                                                                                                                                  
 439   |14900 MHz           |6.8E-01               |+/-.01       |Jy                  |1.49E+10 |6.80E-01    |1.00E-02                  |1.00E-02                  |                           |                           |+/-1.00E-02    |Jy       |1976AJ.....81.1084G|uncertainty                   |14900   MHz        |Broad-band measurement                                                 |024007.09 -001330.7 (B1950)      |Not reported in paper                                   |From Kuhr catalog (1981A&AS...45..367K) |Transformed from previously published data                                                                                                                         
 440   |10.7 GHz (NRAO)     |1.0E+00               |+/-0.03      |Jy                  |1.07E+10 |1.00E+00    |3.00E-02                  |3.00E-02                  |                           |                           |+/-3.00E-02    |Jy       |1973AJ.....78..828K|uncertainty                   |10.7   GHz         |Broad-band measurement                                                 |                                 |Total flux                                              |                                        |From new raw data                                                                                                                                                  
 441   |10695 MHz           |1.0E+00               |+/-.04       |Jy                  |1.07E+10 |1.02E+00    |4.00E-02                  |4.00E-02                  |                           |                           |+/-4.00E-02    |Jy       |1978AJ.....83..451P|uncertainty                   |10695   MHz        |Broad-band measurement                                                 |024007.09 -001330.7 (B1950)      |Not reported in paper                                   |From Kuhr catalog (1981A&AS...45..367K) |Transformed from previously published data                                                                                                                         
 442   |8870 MHz            |1.2E+00               |+/-.05       |Jy                  |8.87E+09 |1.20E+00    |5.00E-02                  |5.00E-02                  |                           |                           |+/-5.00E-02    |Jy       |1973AuJPh..26...93S|uncertainty                   |8870   MHz         |Broad-band measurement                                                 |024007.09 -001330.7 (B1950)      |Not reported in paper                                   |From Kuhr catalog (1981A&AS...45..367K) |Transformed from previously published data                                                                                                                         
 443   |8.46 GHz (VLA)      |9.8E+02               |+/-12.0      |milliJy             |8.46E+09 |9.80E-01    |1.20E-02                  |1.20E-02                  |                           |                           |+/-1.20E-02    |Jy       |2011ApJ...732...45S|rms uncertainty               |8.46 GHz           |Broad-band measurement                                                 |                                 |Total flux                                              |                                        |From new raw data                                                                                                                                                  
 444   |8400 MHz            |1.1E+00               |             |Jy                  |8.40E+09 |1.07E+00    |                          |                          |                           |                           |               |Jy       |1990PKS90.C...0000W|no uncertainty reported       |8400   MHz         |Broad-band measurement                                                 |02 40 07.1 -00 13 31 (B1950)     |Integrated from scans                                   |                                        |Homogenized from new and previously published data                                                                                                                 
 445   |8.4 GHz (VLBA)      |5.4E+00               |+/-0.5       |milliJy             |8.40E+09 |5.40E-03    |5.00E-04                  |5.00E-04                  |                           |                           |+/-5.00E-04    |Jy       |2004ApJ...613..794G|uncertainty                   |8.4 GHz            |Broad-band measurement                                                 |                                 |Flux integrated from map                                |Nuclear flux                            |From new raw data                                                                                                                                                  
 446   |8000 MHz            |1.5E+00               |+/-1.9 %     |Jy                  |8.00E+09 |1.48E+00    |2.81E-02                  |2.81E-02                  |                           |                           |+/-2.81E-02    |Jy       |1971AJ.....76....1S|mean error                    |8000   MHz         |Broad-band measurement                                                 |                                 |Integrated from scans                                   |                                        |From new raw data                                                                                                                                                  
 447   |6.7 GHz (Effelsberg)|1.4E+03               |+/-15  %     |milliJy             |6.70E+09 |1.39E+00    |2.08E-01                  |2.08E-01                  |                           |                           |+/-2.08E-01    |Jy       |2008A&A...484L..43I|estimated error               |6.7 GHz            |Broad-band measurement                                                 |                                 |Flux integrated from map                                |                                        |From new raw data                                                                                                                                                  
 448   |5010 MHz            |1.9E+00               |+/-0.189     |Jy                  |5.01E+09 |1.89E+00    |1.89E-01                  |1.89E-01                  |                           |                           |+/-1.89E-01    |Jy       |1970ApL.....5...29W|estimated error               |5010       MHz     |Broad-band measurement                                                 |                                 |Flux in fixed aperture                                  |                                        |From new raw data                                                                                                                                                  
 449   |5009 MHz            |2.0E+00               |+/-.04       |Jy                  |5.01E+09 |2.01E+00    |4.00E-02                  |4.00E-02                  |                           |                           |+/-4.00E-02    |Jy       |1981A&AS...45..367K|uncertainty                   |5009   MHz         |Broad-band measurement                                                 |024007.09 -001330.7 (B1950)      |Not reported in paper                                   |Recal. to Baars scale by factor of 1.03 |Recalibrated data                                                                                                                                                  
 450   |5009 MHz            |2.0E+00               |+/-.09       |Jy                  |5.01E+09 |1.98E+00    |9.00E-02                  |9.00E-02                  |                           |                           |+/-9.00E-02    |Jy       |1981A&AS...45..367K|uncertainty                   |5009   MHz         |Broad-band measurement                                                 |024007.09 -001330.7 (B1950)      |Not reported in paper                                   |Recal. to Baars scale by factor of 1.03 |Recalibrated data                                                                                                                                                  
 451   |5.0 GHz (VLBA)      |9.1E+00               |+/-0.8       |milliJy             |5.00E+09 |9.10E-03    |8.00E-04                  |8.00E-04                  |                           |                           |+/-8.00E-04    |Jy       |2004ApJ...613..794G|uncertainty                   |5.0 GHz            |Broad-band measurement                                                 |                                 |Flux integrated from map                                |Nuclear flux                            |From new raw data                                                                                                                                                  
 452   |5000 MHz            |1.9E+00               |+/-5   %     |Jy                  |5.00E+09 |1.90E+00    |1.00E-01                  |1.00E-01                  |                           |                           |+/-1.00E-01    |Jy       |1969ApJ...157....1K|rms uncertainty               |5000       MHz     |Broad-band measurement                                                 |                                 |Flux integrated from map                                |                                        |From new raw data                                                                                                                                                  
 453   |5000 MHz            |1.9E+00               |             |Jy                  |5.00E+09 |1.92E+00    |                          |                          |                           |                           |               |Jy       |1990PKS90.C...0000W|no uncertainty reported       |5000   MHz         |Broad-band measurement                                                 |02 40 07.1 -00 13 31 (B1950)     |Integrated from scans                                   |                                        |Homogenized from new and previously published data                                                                                                                 
 454   |5000 MHz            |1.8E+00               |+/-.02       |Jy                  |5.00E+09 |1.83E+00    |2.00E-02                  |2.00E-02                  |                           |                           |+/-2.00E-02    |Jy       |1972AJ.....77..797P|uncertainty                   |5000   MHz         |Broad-band measurement                                                 |024007.09 -001330.7 (B1950)      |Not reported in paper                                   |From Kuhr catalog (1981A&AS...45..367K) |Transformed from previously published data                                                                                                                         
 455   |5000 MHz (NRAO)     |2.2E+00               |+/-0.322     |Jy                  |5.00E+09 |2.19E+00    |3.22E-01                  |3.22E-01                  |                           |                           |+/-3.22E-01    |Jy       |1976ApJS...32..171S|uncertainty                   |5000 MHz           |Broad-band measurement                                                 |02 40 07.7 -00 13 15 (B1950)     |Flux integrated from map                                |                                        |From new raw data                                                                                                                                                  
 456   |5 GHz (VLA)         |1.3E+03               |             |milliJy             |5.00E+09 |1.34E+00    |                          |                          |                           |                           |               |Jy       |2006AJ....132..546G|no uncertainty reported       |5   GHz            |Broad-band measurement                                                 |02 42 40.718 -00 00 46.80 (J2000)|Flux integrated from map                                |Point source flux                       |From new raw data                                                                                                                                                  
 457   |5 GHz (VLA)         |6.6E+02               |             |milliJy             |5.00E+09 |6.64E-01    |                          |                          |                           |                           |               |Jy       |2006AJ....132..546G|no uncertainty reported       |5   GHz            |Broad-band measurement                                                 |02 42 40.718 -00 00 46.80 (J2000)|Flux integrated from map                                |Extranuclear KSR emission; 15" extent   |Averaged from previously published data                                                                                                                            
 458   |5000 MHz            |1.9E+00               |+/-.09       |Jy                  |5.00E+09 |1.89E+00    |9.00E-02                  |9.00E-02                  |                           |                           |+/-9.00E-02    |Jy       |1981A&AS...45..367K|uncertainty                   |5000   MHz         |Broad-band measurement                                                 |024007.09 -001330.7 (B1950)      |Not reported in paper                                   |Recal. to Baars scale by factor of 0.993|Recalibrated data                                                                                                                                                  
 459   |4.89 GHz (VLA)      |1.8E+03               |+/-90        |milliJy             |4.89E+09 |1.80E+00    |9.00E-02                  |9.00E-02                  |                           |                           |+/-9.00E-02    |Jy       |1987ApJ...313..651E|uncertainty                   |4.89   GHz         |Broad-band measurement                                                 |02 40 07.06 -00 13 30.3 (B1950)  |Flux integrated from map                                |Low-resolution data                     |From new raw data                                                                                                                                                  
 460   |4.89 GHz (VLA)      |1.3E+03               |+/-68        |milliJy             |4.89E+09 |1.33E+00    |6.80E-02                  |6.80E-02                  |                           |                           |+/-6.80E-02    |Jy       |1987ApJ...313..651E|uncertainty                   |4.89   GHz         |Broad-band measurement                                                 |02 40 07.06 -00 13 30.3 (B1950)  |Flux integrated from map                                |High-resolution data                    |From new raw data                                                                                                                                                  
 461   |4.86 GHz (VLA)      |1.6E+03               |+/-34.0      |milliJy             |4.86E+09 |1.62E+00    |3.40E-02                  |3.40E-02                  |                           |                           |+/-3.40E-02    |Jy       |2011ApJ...732...45S|rms uncertainty               |4.86 GHz           |Broad-band measurement                                                 |                                 |Total flux                                              |                                        |From new raw data                                                                                                                                                  
 462   |4.85 GHz            |2.0E+03               |+/-99        |milliJy             |4.85E+09 |2.04E+00    |9.90E-02                  |9.90E-02                  |                           |                           |+/-9.90E-02    |Jy       |1995ApJS...97..347G|rms noise                     |4.85       GHz     |Broad-band measurement                                                 |024241.4 -000044 (J2000)         |Modelled datum                                          |                                        |From new raw data; Corrected for contaminating sources                                                                                                             
 463   |4.85 GHz            |2.2E+03               |+/-15  %     |milliJy             |4.85E+09 |2.19E+00    |3.28E-01                  |3.28E-01                  |                           |                           |+/-3.28E-01    |Jy       |1991ApJS...75....1B|uncertainty                   |4.85       GHz     |Broad-band measurement                                                 |024006.9 -001345 (B1950)         |Flux integrated from map                                |                                        |From new raw data; Corrected for contaminating sources                                                                                                             
 464   |4775 MHz (NRAO)     |1.8E+03               |             |milliJy             |4.78E+09 |1.77E+00    |                          |                          |                           |                           |               |Jy       |1986ApJS...61....1B|no uncertainty reported       |4775   MHz         |Broad-band measurement                                                 |02 42 40.4 -00 00 53 (J2000)     |Flux integrated from map                                |S/N = 99.9                              |From new raw data                                                                                                                                                  
 465   |2700 MHz            |3.1E+00               |+/-.15       |Jy                  |2.70E+09 |3.05E+00    |1.50E-01                  |1.50E-01                  |                           |                           |+/-1.50E-01    |Jy       |1981A&AS...45..367K|uncertainty                   |2700   MHz         |Broad-band measurement                                                 |024007.09 -001330.7 (B1950)      |Not reported in paper                                   |Recal. to Baars scale by factor of 1.022|Recalibrated data                                                                                                                                                  
 466   |2700 MHz            |3.3E+00               |             |Jy                  |2.70E+09 |3.27E+00    |                          |                          |                           |                           |               |Jy       |1990PKS90.C...0000W|no uncertainty reported       |2700   MHz         |Broad-band measurement                                                 |02 40 07.1 -00 13 31 (B1950)     |Integrated from scans                                   |                                        |Homogenized from new and previously published data                                                                                                                 
 467   |2700 MHz            |3.1E+00               |+/-.11       |Jy                  |2.70E+09 |3.14E+00    |1.10E-01                  |1.10E-01                  |                           |                           |+/-1.10E-01    |Jy       |1971AuJPA..19....1W|uncertainty                   |2700   MHz         |Broad-band measurement                                                 |024007.09 -001330.7 (B1950)      |Not reported in paper                                   |From Kuhr catalog (1981A&AS...45..367K) |Transformed from previously published data                                                                                                                         
 468   |2700 MHz            |3.2E+00               |+/-.03       |Jy                  |2.70E+09 |3.19E+00    |3.00E-02                  |3.00E-02                  |                           |                           |+/-3.00E-02    |Jy       |1975AuJPA..38....1W|uncertainty                   |2700   MHz         |Broad-band measurement                                                 |024007.09 -001330.7 (B1950)      |Not reported in paper                                   |From Kuhr catalog (1981A&AS...45..367K) |Transformed from previously published data                                                                                                                         
 469   |2695 MHz            |3.0E+00               |+/-.05       |Jy                  |2.70E+09 |3.02E+00    |5.00E-02                  |5.00E-02                  |                           |                           |+/-5.00E-02    |Jy       |1981A&AS...45..367K|uncertainty                   |2695   MHz         |Broad-band measurement                                                 |024007.09 -001330.7 (B1950)      |Not reported in paper                                   |Recal. to Baars scale by factor of 1.011|Recalibrated data                                                                                                                                                  
 470   |2695 MHz            |2.8E+00               |+/-.22       |Jy                  |2.70E+09 |2.80E+00    |2.20E-01                  |2.20E-01                  |                           |                           |+/-2.20E-01    |Jy       |1972MNRAS.159..233A|uncertainty                   |2695   MHz         |Broad-band measurement                                                 |024007.09 -001330.7 (B1950)      |Not reported in paper                                   |From Kuhr catalog (1981A&AS...45..367K) |Transformed from previously published data                                                                                                                         
 471   |2695 MHz            |3.0E+00               |+/-5   %     |Jy                  |2.70E+09 |2.99E+00    |1.50E-01                  |1.50E-01                  |                           |                           |+/-1.50E-01    |Jy       |1969ApJ...157....1K|rms uncertainty               |2695       MHz     |Broad-band measurement                                                 |                                 |Flux integrated from map                                |                                        |From new raw data                                                                                                                                                  
 472   |2650 MHz            |3.2E+00               |+/-.03       |Jy                  |2.65E+09 |3.18E+00    |3.00E-02                  |3.00E-02                  |                           |                           |+/-3.00E-02    |Jy       |1975AuJPA..38....1W|uncertainty                   |2650   MHz         |Broad-band measurement                                                 |024007.09 -001330.7 (B1950)      |Not reported in paper                                   |From Kuhr catalog (1981A&AS...45..367K) |Transformed from previously published data                                                                                                                         
 473   |1465 MHz            |5.0E+03               |+/-230       |milliJy             |1.46E+09 |4.96E+00    |2.30E-01                  |2.30E-01                  |                           |                           |+/-2.30E-01    |Jy       |1983ApJS...53..459C|rms uncertainty               |1465       MHz     |Broad-band measurement                                                 |                                 |Flux integrated from map                                |                                        |From new raw data                                                                                                                                                  
 474   |1.46 GHz (VLA)      |4.6E+03               |+/-230       |milliJy             |1.46E+09 |4.61E+00    |2.30E-01                  |2.30E-01                  |                           |                           |+/-2.30E-01    |Jy       |1987ApJ...313..651E|uncertainty                   |1.46   GHz         |Broad-band measurement                                                 |02 40 07.06 -00 13 30.3 (B1950)  |Flux integrated from map                                |                                        |From new raw data                                                                                                                                                  
 483   |1410 MHz            |5.4E+00               |+/-.13       |Jy                  |1.41E+09 |5.44E+00    |1.30E-01                  |1.30E-01                  |                           |                           |+/-1.30E-01    |Jy       |1981A&AS...45..367K|uncertainty                   |1410   MHz         |Broad-band measurement                                                 |024007.09 -001330.7 (B1950)      |Not reported in paper                                   |Recal. to Baars scale by factor of 1.017|Recalibrated data                                                                                                                                                  
 484   |1410 MHz            |5.1E+00               |             |Jy                  |1.41E+09 |5.10E+00    |                          |                          |                           |                           |               |Jy       |1990PKS90.C...0000W|no uncertainty reported       |1410   MHz         |Broad-band measurement                                                 |02 40 07.1 -00 13 31 (B1950)     |Integrated from scans                                   |                                        |Homogenized from new and previously published data                                                                                                                 
 485   |1.4 GHz (VLA)       |4.9E+03               |             |milliJy             |1.40E+09 |4.85E+00    |                          |                          |                           |                           |               |Jy       |2002AJ....124..675C|no uncertainty reported       |1.4   GHz          |Broad-band measurement                                                 |                                 |Flux integrated from map                                |                                        |Averaged from previously published data                                                                                                                            
 486   |1.4 GHz (VLBA)      |                      |<0.06        |milliJy             |1.40E+09 |            |                          |                          |0.00006000                 |                           |<6.00E-05      |Jy       |2004ApJ...613..794G|uncertainty                   |1.4 GHz            |Broad-band measurement                                                 |                                 |Flux integrated from map                                |Nuclear flux                            |From new raw data                                                                                                                                                  
 487   |1400 MHz            |5.0E+00               |+/-.14       |Jy                  |1.40E+09 |5.04E+00    |1.40E-01                  |1.40E-01                  |                           |                           |+/-1.40E-01    |Jy       |1981A&AS...45..367K|uncertainty                   |1400   MHz         |Broad-band measurement                                                 |024007.09 -001330.7 (B1950)      |Not reported in paper                                   |Recal. to Baars scale by factor of 1.029|Recalibrated data                                                                                                                                                  
 488   |1400 MHz            |4.9E+00               |+/-5   %     |Jy                  |1.40E+09 |4.90E+00    |2.40E-01                  |2.40E-01                  |                           |                           |+/-2.40E-01    |Jy       |1969ApJ...157....1K|rms uncertainty               |1400       MHz     |Broad-band measurement                                                 |                                 |Flux integrated from map                                |                                        |From new raw data                                                                                                                                                  
 489   |1.40 GHz            |4.8E+03               |             |milliJy             |1.40E+09 |4.85E+00    |                          |                          |                           |                           |               |Jy       |1992ApJS...79..331W|no uncertainty reported       |1.4        GHz     |Broad-band measurement                                                 |024006.9 -001345 (B1950)         |Peak flux                                               |                                        |From new raw data                                                                                                                                                  
 490   |1400 MHz            |5.0E+00               |+/-.30       |Jy                  |1.40E+09 |5.00E+00    |3.00E-01                  |3.00E-01                  |                           |                           |+/-3.00E-01    |Jy       |1981A&AS...45..367K|uncertainty                   |1400   MHz         |Broad-band measurement                                                 |024007.09 -001330.7 (B1950)      |Not reported in paper                                   |Recal. to Baars scale by factor of 1.029|Recalibrated data                                                                                                                                                  
 491   |1400 MHz (NRAO)     |5.0E+00               |+/-0.09      |Jy                  |1.40E+09 |4.97E+00    |9.00E-02                  |9.00E-02                  |                           |                           |+/-9.00E-02    |Jy       |1966ApJS...13...65P|internal error                |1400       MHz     |Broad-band measurement                                                 |024006.3 -001337. (B1950)        |Peak flux                                               |                                        |From new raw data                                                                                                                                                  
 492   |1400 MHz (NRAO)     |4.9E+00               |             |Jy                  |1.40E+09 |4.90E+00    |                          |                          |                           |                           |               |Jy       |1964AJ.....69..277H|no uncertainty reported       |1400      MHz      |Broad-band measurement; peak value reported                            |024007 -0014 (B1950)             |Peak flux                                               |                                        |From new raw data                                                                                                                                                  
 493   |960 MHz             |6.8E+00               |+/-.13       |Jy                  |9.60E+08 |6.82E+00    |1.30E-01                  |1.30E-01                  |                           |                           |+/-1.30E-01    |Jy       |1981A&AS...45..367K|uncertainty                   |960   MHz          |Broad-band measurement                                                 |024007.09 -001330.7 (B1950)      |Not reported in paper                                   |Recal. to Baars scale by factor of 1.029|Recalibrated data                                                                                                                                                  
 494   |750 MHz (NRAO)      |7.5E+00               |             |Jy                  |7.50E+08 |7.50E+00    |                          |                          |                           |                           |               |Jy       |1964AJ.....69..277H|no uncertainty reported       |750      MHz       |Broad-band measurement; peak value reported                            |024007 -0014 (B1950)             |Peak flux                                               |                                        |From new raw data                                                                                                                                                  
 495   |750 MHz             |7.6E+00               |+/-.40       |Jy                  |7.50E+08 |7.60E+00    |4.00E-01                  |4.00E-01                  |                           |                           |+/-4.00E-01    |Jy       |1981A&AS...45..367K|uncertainty                   |750   MHz          |Broad-band measurement                                                 |024007.09 -001330.7 (B1950)      |Not reported in paper                                   |Recal. to Baars scale by factor of 1.046|Recalibrated data                                                                                                                                                  
 496   |750 MHz             |7.3E+00               |+/-5   %     |Jy                  |7.50E+08 |7.30E+00    |3.60E-01                  |3.60E-01                  |                           |                           |+/-3.60E-01    |Jy       |1969ApJ...157....1K|rms uncertainty               |750        MHz     |Broad-band measurement                                                 |                                 |Flux integrated from map                                |                                        |From new raw data                                                                                                                                                  
 497   |750 MHz             |8.1E+00               |+/-.11       |Jy                  |7.50E+08 |8.09E+00    |1.10E-01                  |1.10E-01                  |                           |                           |+/-1.10E-01    |Jy       |1981A&AS...45..367K|uncertainty                   |750   MHz          |Broad-band measurement                                                 |024007.09 -001330.7 (B1950)      |Not reported in paper                                   |Recal. to Baars scale by factor of 1.059|Recalibrated data                                                                                                                                                  
 498   |750 MHz (NRAO)      |7.6E+00               |+/-0.10      |Jy                  |7.50E+08 |7.64E+00    |1.00E-01                  |1.00E-01                  |                           |                           |+/-1.00E-01    |Jy       |1966ApJS...13...65P|internal error                |750        MHz     |Broad-band measurement                                                 |024006.3 -001337. (B1950)        |Peak flux                                               |                                        |From new raw data                                                                                                                                                  
 499   |635 MHz             |9.4E+00               |+/-.28       |Jy                  |6.35E+08 |9.43E+00    |2.80E-01                  |2.80E-01                  |                           |                           |+/-2.80E-01    |Jy       |1981A&AS...45..367K|uncertainty                   |635   MHz          |Broad-band measurement                                                 |024007.09 -001330.7 (B1950)      |Not reported in paper                                   |Recal. to Baars scale by factor of 1.035|Recalibrated data                                                                                                                                                  
 500   |635 MHz             |8.5E+00               |             |Jy                  |6.35E+08 |8.50E+00    |                          |                          |                           |                           |               |Jy       |1990PKS90.C...0000W|no uncertainty reported       |635   MHz          |Broad-band measurement                                                 |02 40 07.1 -00 13 31 (B1950)     |Integrated from scans                                   |                                        |Homogenized from new and previously published data                                                                                                                 
 501   |468 MHz             |1.1E+01               |+/-.85       |Jy                  |4.68E+08 |1.12E+01    |8.50E-01                  |8.50E-01                  |                           |                           |+/-8.50E-01    |Jy       |1981A&AS...45..367K|uncertainty                   |468   MHz          |Broad-band measurement                                                 |024007.09 -001330.7 (B1950)      |Not reported in paper                                   |Recal. to Baars scale by factor of 1.045|Recalibrated data                                                                                                                                                  
 502   |408 MHz             |1.2E+01               |             |Jy                  |4.08E+08 |1.24E+01    |                          |                          |                           |                           |               |Jy       |1990PKS90.C...0000W|no uncertainty reported       |408   MHz          |Broad-band measurement                                                 |02 40 07.1 -00 13 31 (B1950)     |Integrated from scans                                   |                                        |Homogenized from new and previously published data                                                                                                                 
 503   |408 MHz             |1.2E+01               |+/-0.54      |Jy                  |4.08E+08 |1.24E+01    |5.40E-01                  |5.40E-01                  |                           |                           |+/-5.40E-01    |Jy       |1981MNRAS.194..693L|rms noise                     |408        MHz     |Broad-band measurement                                                 |024007.1 -001321 (B1950)         |Modelled datum                                          |                                        |From new raw data; Corrected for contaminating sources                                                                                                             
 504   |408 MHz             |1.0E+01               |+/-2.52      |Jy                  |4.08E+08 |1.01E+01    |2.52E+00                  |2.52E+00                  |                           |                           |+/-2.52E+00    |Jy       |1969AuJPA...7....3E|uncertainty                   |408   MHz          |Broad-band measurement                                                 |024007.09 -001330.7 (B1950)      |Not reported in paper                                   |From Kuhr catalog (1981A&AS...45..367K) |Transformed from previously published data                                                                                                                         
 505   |365 MHz (Texas)     |1.1E+01               |+/-0.179     |Jy                  |3.65E+08 |1.14E+01    |1.79E-01                  |1.79E-01                  |                           |                           |+/-1.79E-01    |Jy       |1996AJ....111.1945D|internal error                |365        MHz     |Broad-band measurement; obtained by interpolation over frequency       |024007.064 -001330.93 (B1950)    |Integrated from scans                                   |Model:D;MFlag:+;EFlag:+;LFlag:+.        |From new raw data                                                                                                                                                  
 506   |318 MHz             |1.2E+01               |+/-.49       |Jy                  |3.18E+08 |1.23E+01    |4.90E-01                  |4.90E-01                  |                           |                           |+/-4.90E-01    |Jy       |1981A&AS...45..367K|uncertainty                   |318   MHz          |Broad-band measurement                                                 |024007.09 -001330.7 (B1950)      |Not reported in paper                                   |Recal. to Baars scale by factor of 1.05 |Recalibrated data                                                                                                                                                  
 507   |178 MHz             |1.6E+01               |+/-15  %     |Jy                  |1.78E+08 |1.61E+01    |2.42E+00                  |2.42E+00                  |                           |                           |+/-2.42E+00    |Jy       |1969ApJ...157....1K|rms uncertainty               |178        MHz     |Broad-band measurement                                                 |                                 |Flux integrated from map                                |                                        |From new raw data                                                                                                                                                  
 508   |178 MHz             |1.7E+01               |+/-1.70      |Jy                  |1.78E+08 |1.73E+01    |1.70E+00                  |1.70E+00                  |                           |                           |+/-1.70E+00    |Jy       |1981A&AS...45..367K|uncertainty                   |178   MHz          |Broad-band measurement                                                 |024007.09 -001330.7 (B1950)      |Not reported in paper                                   |Recal. to Baars scale by factor of 1.19 |Recalibrated data                                                                                                                                                  
 509   |178 MHz             |1.8E+01               |+/-1.80      |Jy                  |1.78E+08 |1.79E+01    |1.80E+00                  |1.80E+00                  |                           |                           |+/-1.80E+00    |Jy       |1981A&AS...45..367K|uncertainty                   |178   MHz          |Broad-band measurement                                                 |024007.09 -001330.7 (B1950)      |Not reported in paper                                   |Recal. to Baars scale by factor of 1.11 |Recalibrated data                                                                                                                                                  
 510   |178 MHz             |1.6E+01               |+/-8.0 %     |Jy                  |1.78E+08 |1.61E+01    |1.29E+00                  |1.29E+00                  |                           |                           |+/-1.29E+00    |Jy       |1967MmRAS..71...49G|uncertainty                   |178        MHz     |Broad-band measurement                                                 |024005.9 -001300 (B1950)         |Integrated from scans                                   |                                        |From new raw data; Uncorrected for known sources in beam                                                                                                           
 511   |178 MHz             |1.6E+01               |             |Jy                  |1.78E+08 |1.61E+01    |                          |                          |                           |                           |               |Jy       |1990PKS90.C...0000W|no uncertainty reported       |178   MHz          |Broad-band measurement                                                 |02 40 07.1 -00 13 31 (B1950)     |Integrated from scans                                   |                                        |Homogenized from new and previously published data                                                                                                                 
 512   |160 MHz             |2.1E+01               |             |Jy                  |1.60E+08 |2.05E+01    |                          |                          |                           |                           |               |Jy       |1995AuJPh..48..143S|no uncertainty reported       |160        MHz     |Broad-band measurement                                                 |024007.8 -001217. (B1950)        |Flux integrated from map                                |                                        |From new raw data                                                                                                                                                  
 513   |160 MHz             |2.1E+01               |+/-3.20      |Jy                  |1.60E+08 |2.14E+01    |3.20E+00                  |3.20E+00                  |                           |                           |+/-3.20E+00    |Jy       |1981A&AS...45..367K|uncertainty                   |160   MHz          |Broad-band measurement                                                 |024007.09 -001330.7 (B1950)      |Not reported in paper                                   |Recal. to Baars scale by factor of 1.11 |Recalibrated data                                                                                                                                                  
 514   |145 MHz (PAPER)     |2.1E+01               |             |Jy                  |1.45E+08 |2.14E+01    |                          |                          |                           |                           |               |Jy       |2011ApJ...734L..34J|no uncertainty reported       |145 MHz            |Broad-band measurement                                                 |40.87 0.15 (J2000)               |Flux integrated from map                                |                                        |From new raw data                                                                                                                                                  
 515   |80 MHz              |2.4E+01               |             |Jy                  |8.00E+07 |2.40E+01    |                          |                          |                           |                           |               |Jy       |1995AuJPh..48..143S|no uncertainty reported       |80        MHz      |Broad-band measurement                                                 |024007.8 -001217. (B1950)        |Flux integrated from map                                |                                        |From new raw data                                                                                                                                                  
 516   |80 MHz              |2.2E+01               |             |Jy                  |8.00E+07 |2.20E+01    |                          |                          |                           |                           |               |Jy       |1990PKS90.C...0000W|no uncertainty reported       |80   MHz           |Broad-band measurement                                                 |02 40 07.1 -00 13 31 (B1950)     |Integrated from scans                                   |                                        |Homogenized from new and previously published data                                                                                                                 
 517   |80 MHz              |2.4E+01               |+/-4.00      |Jy                  |8.00E+07 |2.40E+01    |4.00E+00                  |4.00E+00                  |                           |                           |+/-4.00E+00    |Jy       |1981A&AS...45..367K|uncertainty                   |80   MHz           |Broad-band measurement                                                 |024007.09 -001330.7 (B1950)      |Not reported in paper                                   |Recal. to Baars scale by factor of 1.074|Recalibrated data                                                                                                                                                  
 518   |74 MHz (VLA)        |2.7E+01               |+/-2.80      |Jy                  |7.38E+07 |2.73E+01    |2.80E+00                  |2.80E+00                  |                           |                           |+/-2.80E+00    |Jy       |2007AJ....134.1245C|rms uncertainty               |73.8   MHz         |Broad-band measurement                                                 |02 42 40.84 -00 00 45.4 (J2000)  |Flux integrated from map                                |Corrected for clean bias                |From new raw data                                                                                                                                                  
 519   |57.5 MHz            |3.9E+01               |+/-8.0       |Jy                  |5.75E+07 |3.90E+01    |8.00E+00                  |8.00E+00                  |                           |                           |+/-8.00E+00    |Jy       |1990ApJ...352...30I|uncertainty                   |57.5       MHz     |Broad-band measurement                                                 |                                 |Flux integrated from map                                |                                        |From new raw data                                                                                                                                                  
 520   |38 MHz              |3.3E+01               |+/-25  %     |Jy                  |3.80E+07 |3.30E+01    |8.25E+00                  |8.25E+00                  |                           |                           |+/-8.25E+00    |Jy       |1969ApJ...157....1K|rms uncertainty               |38         MHz     |Broad-band measurement                                                 |                                 |Flux integrated from map                                |                                        |From new raw data                                                                                                                                                  
 521   |22 MHz (DRAO)       |8.3E+01               |+/-8         |Jy                  |2.23E+07 |8.30E+01    |8.00E+00                  |8.00E+00                  |                           |                           |+/-8.00E+00    |Jy       |1986A&AS...65..485R|uncertainty                   |22.25 MHz          |Broad-band measurement                                                 |02 40 06.0 -00 25 00 (B1950)     |Flux integrated from map                                |                                        |From new raw data                                                                                                                                                  
