
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-02-19T10:33:25PST



Photometric Data for ERO N4

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
4|16 microns (Spitzer/IRS)| 0.52      |+/-10  %| milliJy            |1.86E+13|  5.20E-04|+/-5.20E-05|Jy|2004ApJS..154..142C|uncertainty|     16.10 microns   | Broad-band measurement|04 43 07.1 +02 10 25.1 (J2000)| Flux integrated from map|                                        |From new raw data
5|22 microns (Spitzer/IRS)| 0.98      |+/-10  %| milliJy            |1.35E+13|  9.80E-04|+/-9.80E-05|Jy|2004ApJS..154..142C|uncertainty|     22.25 microns   | Broad-band measurement|04 43 07.1 +02 10 25.1 (J2000)| Flux integrated from map|                                        |From new raw data
7|450 microns (SCUBA) | |<60        |milliJy             |6.66E+11| |6.00E-02|Jy|2002MNRAS.331..495S|3rms uncertainty reported|     450   microns   | Broad-band measurement|044307.2 +021024 (J2000)| Flux integrated from map|                                        |From new raw data
8|850 microns (SCUBA) | 7.2       |1.5 |milliJy             |3.53E+11|  7.20E-03|1.50E-03 |Jy|2002MNRAS.331..495S|no uncertainty reported|     850   microns   | Broad-band measurement|044307.2 +021024 (J2000)| Flux integrated from map|                                        |From new raw data
10|1.3 mm (PdBI)      | |<1.2       |milliJy             |2.31E+11| |1.20E-03|Jy|2006ApJ...640..228T|3rms uncertainty reported|     1.3   mm        | Broad-band measurement| | Flux integrated from map|                                        |From new raw data
