
Results from query to  NASA/IPAC Extragalactic Database (NED),
which is operated by the Jet Propulsion Laboratory, California Institute of
Technology, under contract with the National Aeronautics and Space Administration.
This work was (partially) supported by the US National Virtual Observatory
development project, which is funded by the National Science Foundation
under cooperative agreement AST0122449 with The Johns Hopkins University.



queryDateTime:2013-05-28T01:42:09PDT



Photometric Data for SPT-S053816-5030.8, z=2.783

No.|Observed Passband|Photometry Measurement|Uncertainty|Units|Frequency|NED Photometry Measurement|NED Uncertainty|NED Units|Refcode|Significance|Published frequency|Frequency Mode|Coordinates Targeted|Spatial Mode|Qualifiers|Comments
1|3.6 microns (IRAC) | 0.022     |+/-0.005|mJy             |8.44E+13|  0.022E-03|+/-0.005E-03|Jy|2011ApJ...728L...4H|uncertainty|     3.550 microns   | Broad-band measurement|09 13 05.0 -00 53 43 (J2000)| Flux in fixed aperture|                                        |From new raw data
2|4.5 microns (IRAC) | 0.047     |+/-0.008|mJy             |6.67E+13|  0.047E-03|+/-0.008E-03|Jy|2011ApJ...728L...4H|uncertainty|     4.493 microns   | Broad-band measurement|09 13 05.0 -00 53 43 (J2000)| Flux in fixed aperture|                                        |From new raw data
3|100 microns (PACS) | 31.       |+/-2.0  |mJy             |2.998e+12| 31.E-03 |+/-2.0E-03|Jy|2005MNRAS.358..149P|1rms uncertainty|     850   microns   | Broad-band measurement|12 37 11.7 +62 22 12 (J2000)| Flux integrated from map|                                        |Averaged new and previously published data
4|160 microns (PACS) | 141.0     |+/-15.0 |mJy             |1.874e+12| 141.E-03|+/-15.0E-03 |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
5|250 microns (SPIRE)| 326.      |+/-23.0 |mJy             |1.199e+12| 326.0E-03|+/-23.0e-03 |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
6|350 microns (SPIRE)| 396.      |+/-38.  |mJy             |8.565e+11|396.E-03 |+/-38.0e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
7|352 microns (APEX) | 336.      |+/-88.  |mJy             |8.52E+11|  336.0E-03|+/-88.0E-03|Jy|2010Natur.464..733S|uncertainty|       352 microns   | Broad-band measurement|21 35 11.6 -01 02 52.0 (J2000)| Flux in fixed aperture|                                        |From new raw data
8|500 microns (SPIRE) | 325.     |+/-24.0 |mJy             |5.996e+11|325.E-03 |+/-24.0e-03  |Jy |2.40e+01 |0.00e+00 |-9.90e+01 |-9.90e+01 |-9.90e+01 | NaN|
9|870 microns (APEX) | 125       |+/-7    |mJy             |3.45E+11|  125.0E-03|+/-7.0E-03 |Jy|2010Natur.464..733S|uncertainty|       870 microns   | Broad-band measurement|21 35 11.6 -01 02 52.0 (J2000)| Flux in fixed aperture|                                        |From new raw data
10|890 microns (SMA)  | 132.0     |+/-26.4 |mJy             |3.37E+11| 132.0E-3 |+/-26.4E-3 |Jy|2007MNRAS.376.1073Z|no uncertainty reported|     850   microns   | Broad-band measurement|02 39 51.9 -01 35 55 (J2000)| Flux integrated from map|S/N = 19.9                              |From reprocessed raw data
11|1.4mm (SPT) | 28.0      |+/-4.6  |mJy             |2.20436E+11| 28.0E-3|+/-4.6E-3 |Jy|2007MNRAS.376.1073Z|no uncertainty reported|     850   microns   | Broad-band measurement|02 39 51.9 -01 35 55 (J2000)| Flux integrated from map|S/N = 19.9                              |From reprocessed raw data
1|1.4 mm (SPT)        | 31.31     ||milliJy             |2.20E+11|  3.13E-02||Jy|2010ApJ...719..763V|no uncertainty reported|       1.4 mm        | Broad-band measurement|84.569 -50.514 (J2000)| Flux integrated from map|Raw flux; S/N = 9.04                    |From new raw data
2|1.4 mm (SPT)        | 29.68     |+/-4.52 |milliJy             |2.20E+11|  2.97E-02|+/-4.52E-03|Jy|2010ApJ...719..763V|uncertainty|       1.4 mm        | Broad-band measurement|84.569 -50.514 (J2000)| Flux integrated from map|De-boosted flux; S/N = 9.04             |From new raw data
12|2.0mm (SPT) | 8.5       |+/-1.4  |mJy             |1.53740E+11| 8.5E-3 |+/-1.4E-3 |Jy|2007MNRAS.376.1073Z|no uncertainty reported|     850   microns   | Broad-band measurement|02 39 51.9 -01 35 55 (J2000)| Flux integrated from map|S/N = 19.9                              |From reprocessed raw data
3|2.0 mm (SPT)        | 8.54      |+/-1.35 |milliJy             |1.50E+11|  8.54E-03|+/-1.35E-03|Jy|2010ApJ...719..763V|uncertainty|       2.0 mm        | Broad-band measurement|84.569 -50.514 (J2000)| Flux integrated from map|De-boosted flux; S/N = 6.81             |From new raw data
4|2.0 mm (SPT)        | 8.78      ||milliJy             |1.50E+11|  8.78E-03||Jy|2010ApJ...719..763V|no uncertainty reported|       2.0 mm        | Broad-band measurement|84.569 -50.514 (J2000)| Flux integrated from map|Raw flux; S/N = 6.81                    |From new raw data
13|8.6mm (ATCA)       | 0.13      |+/-0.02 |mJy             |3.48596e+10| 0.13E-03|+/-0.02E-03|Jy|2010A&A...518L..35I|3rms uncertainty|      4.49 cm        | Broad-band measurement| | Flux integrated from map|                                        |From new raw data
14|0.85cm (VLA)       |           |<120|microJy             |35.0E+09| |120.0E-06|Jy|2010A&A...518L..35I|3rms uncertainty|      4.49 cm        | Broad-band measurement| | Flux integrated from map|                                        |From new raw data
15|0.97cm (VLA)       |           |<120|microJy             |31.0E+09| |120.0E-06|Jy|2010A&A...518L..35I|3rms uncertainty|      4.49 cm        | Broad-band measurement| | Flux integrated from map|                                        |From new raw data
